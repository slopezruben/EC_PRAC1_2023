//: version "1.8.7"

module CSA(A, Cin, Cout, B, S);
//: interface  /sz:(139, 87) /bd:[ Ti0>B[3:0](94/139) Ti1>A[3:0](41/139) Ri0>Cin(39/87) Lo0<Cout(49/87) Bo0<S[3:0](66/139) ]
input [3:0] B;    //: /sn:0 /dp:1 {0}(508,86)(480,86){1}
//: {2}(479,86)(376,86){3}
//: {4}(375,86)(279,86){5}
//: {6}(278,86)(176,86){7}
//: {8}(175,86)(123,86){9}
input [3:0] A;    //: /sn:0 {0}(468,55)(452,55){1}
//: {2}(451,55)(343,55){3}
//: {4}(342,55)(245,55){5}
//: {6}(244,55)(154,55){7}
//: {8}(153,55)(132,55){9}
input Cin;    //: /sn:0 /dp:17 {0}(437,349)(420,349)(420,369)(387,369)(387,395)(338,395)(338,352){1}
//: {2}(340,350)(352,350){3}
//: {4}(336,350)(228,350)(228,352){5}
//: {6}(230,354)(252,354){7}
//: {8}(226,354)(133,354)(133,355){9}
//: {10}(135,357)(152,357){11}
//: {12}(131,357)(62,357)(62,358)(54,358){13}
//: {14}(52,356)(52,233){15}
//: {16}(52,360)(52,404)(37,404){17}
output Cout;    //: /sn:0 {0}(28,111)(18,111)(18,195)(29,195)(29,210)(39,210){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(310,447)(310,475)(321,475)(321,481)(262,481)(262,495)(321,495){1}
wire w6;    //: /sn:0 {0}(460,362)(460,403)(295,403)(295,441){1}
wire w16;    //: /sn:0 /dp:1 {0}(68,220)(139,220)(139,274)(149,274){1}
wire w7;    //: /sn:0 {0}(391,164)(427,164)(427,166)(437,166){1}
wire w25;    //: /sn:0 {0}(350,270)(325,270)(325,263)(315,263){1}
wire w4;    //: /sn:0 {0}(557,188)(557,161)(500,161){1}
wire w3;    //: /sn:0 {0}(501,244)(501,122)(482,122){1}
//: {2}(480,120)(480,90){3}
//: {4}(480,124)(480,141){5}
wire w22;    //: /sn:0 {0}(392,246)(392,123)(379,123){1}
//: {2}(377,121)(377,96)(376,96)(376,90){3}
//: {4}(377,125)(377,146){5}
wire w0;    //: /sn:0 /dp:1 {0}(450,333)(450,200)(469,200)(469,190){1}
wire w20;    //: /sn:0 {0}(456,268)(421,268)(421,264)(411,264){1}
wire w30;    //: /sn:0 {0}(254,269)(228,269)(228,267)(218,267){1}
wire w29;    //: /sn:0 {0}(275,367)(275,425)(315,425)(315,441){1}
wire w12;    //: /sn:0 {0}(298,167)(320,167)(320,166)(330,166){1}
wire w19;    //: /sn:0 {0}(163,194)(163,332)(165,332)(165,341){1}
wire w18;    //: /sn:0 /dp:1 {0}(265,338)(265,201)(263,201)(263,191){1}
wire w23;    //: /sn:0 {0}(367,246)(367,129)(349,129){1}
//: {2}(347,127)(347,65)(343,65)(343,59){3}
//: {4}(347,131)(347,146){5}
wire w10;    //: /sn:0 {0}(556,285)(556,267)(517,267){1}
wire w21;    //: /sn:0 /dp:1 {0}(285,338)(285,297)(280,297)(280,287){1}
wire w1;    //: /sn:0 /dp:1 {0}(470,333)(470,296)(482,296)(482,286){1}
wire w31;    //: /sn:0 {0}(175,370)(175,385)(325,385)(325,441){1}
wire w32;    //: /sn:0 {0}(196,246)(196,140)(181,140){1}
//: {2}(179,138)(179,96)(176,96)(176,90){3}
//: {4}(179,142)(179,151){5}
wire w8;    //: /sn:0 {0}(473,244)(473,126)(456,126){1}
//: {2}(454,124)(454,65)(452,65)(452,59){3}
//: {4}(454,128)(454,141){5}
wire w17;    //: /sn:0 {0}(198,169)(227,169)(227,173)(237,173){1}
wire w27;    //: /sn:0 {0}(296,245)(296,131)(281,131){1}
//: {2}(279,129)(279,90){3}
//: {4}(279,133)(279,149){5}
wire w28;    //: /sn:0 {0}(271,245)(271,129)(256,129){1}
//: {2}(254,127)(254,65)(245,65)(245,59){3}
//: {4}(254,131)(254,149){5}
wire w33;    //: /sn:0 {0}(168,246)(168,134)(156,134){1}
//: {2}(154,132)(154,59){3}
//: {4}(154,136)(154,151){5}
wire w11;    //: /sn:0 {0}(375,363)(375,415)(305,415)(305,441){1}
wire w15;    //: /sn:0 /dp:1 {0}(68,200)(127,200)(127,175)(137,175){1}
wire w5;    //: /sn:0 /dp:1 {0}(185,341)(185,306)(178,306)(178,296){1}
wire w9;    //: /sn:0 {0}(356,188)(356,324)(365,324)(365,334){1}
wire w26;    //: /sn:0 {0}(376,288)(376,324)(385,324)(385,334){1}
//: enddecls

  FA g4 (.A(w8), .B(w3), .Cin(w10), .Cout(w20), .S(w1));   //: @(457, 245) /sz:(59, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: input g8 (A) @(130,55) /sn:0 /w:[ 9 ]
  FA g3 (.A(w33), .B(w32), .Cin(w17), .Cout(w15), .S(w19));   //: @(138, 152) /sz:(59, 41) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Lo0<1 Bo0<0 ]
  tran g16(.Z(w28), .I(A[2]));   //: @(245,53) /sn:0 /R:1 /w:[ 3 6 5 ] /ss:1
  tran g17(.Z(w33), .I(A[3]));   //: @(154,53) /sn:0 /R:1 /w:[ 3 8 7 ] /ss:1
  //: input g26 (Cin) @(35,404) /sn:0 /w:[ 17 ]
  FA g2 (.A(w28), .B(w27), .Cin(w12), .Cout(w17), .S(w18));   //: @(238, 150) /sz:(59, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Lo0<1 Bo0<1 ]
  //: joint g23 (w23) @(347, 129) /w:[ 1 2 -1 4 ]
  //: output g30 (Cout) @(25,111) /sn:0 /w:[ 0 ]
  FA g1 (.A(w23), .B(w22), .Cin(w7), .Cout(w12), .S(w9));   //: @(331, 147) /sz:(59, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Lo0<1 Bo0<0 ]
  //: joint g24 (w8) @(454, 126) /w:[ 1 2 -1 4 ]
  //: switch g39 (w4) @(557,202) /sn:0 /R:1 /w:[ 0 ] /st:0
  mux g29 (.I0(w15), .I1(w16), .S(Cin), .Z(Cout));   //: @(52,210) /sn:0 /R:3 /delay:" 3 3" /w:[ 0 0 15 1 ] /ss:1 /do:0
  //: joint g18 (w32) @(179, 140) /w:[ 1 2 -1 4 ]
  tran g10(.Z(w3), .I(B[0]));   //: @(480,84) /sn:0 /R:1 /w:[ 3 2 1 ] /ss:1
  //: joint g25 (w3) @(480, 122) /w:[ 1 2 -1 4 ]
  FA g6 (.A(w28), .B(w27), .Cin(w25), .Cout(w30), .S(w21));   //: @(255, 246) /sz:(59, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  FA g7 (.A(w33), .B(w32), .Cin(w30), .Cout(w16), .S(w5));   //: @(150, 247) /sz:(67, 48) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 ]
  //: input g9 (B) @(121,86) /sn:0 /w:[ 9 ]
  //: joint g35 (Cin) @(228, 354) /w:[ 6 5 8 -1 ]
  //: joint g22 (w22) @(377, 123) /w:[ 1 2 -1 4 ]
  mux g31 (.I0(w18), .I1(w21), .S(Cin), .Z(w29));   //: @(275,354) /sn:0 /delay:" 3 3" /w:[ 0 0 7 0 ] /ss:0 /do:0
  //: joint g33 (Cin) @(52, 358) /w:[ 13 14 -1 16 ]
  //: joint g36 (Cin) @(338, 350) /w:[ 2 -1 4 1 ]
  //: switch g40 (w10) @(556,299) /sn:0 /R:1 /w:[ 0 ] /st:1
  tran g12(.Z(w27), .I(B[2]));   //: @(279,84) /sn:0 /R:1 /w:[ 3 6 5 ] /ss:1
  mux g28 (.I0(w9), .I1(w26), .S(Cin), .Z(w11));   //: @(375,350) /sn:0 /delay:" 3 3" /w:[ 1 1 3 0 ] /ss:0 /do:0
  //: joint g34 (Cin) @(133, 357) /w:[ 10 9 12 -1 ]
  FA g5 (.A(w23), .B(w22), .Cin(w20), .Cout(w25), .S(w26));   //: @(351, 247) /sz:(59, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  tran g11(.Z(w22), .I(B[1]));   //: @(376,84) /sn:0 /R:1 /w:[ 3 4 3 ] /ss:1
  tran g14(.Z(w8), .I(A[0]));   //: @(452,53) /sn:0 /R:1 /w:[ 3 2 1 ] /ss:1
  //: joint g19 (w33) @(154, 134) /w:[ 1 2 -1 4 ]
  //: joint g21 (w27) @(279, 131) /w:[ 1 2 -1 4 ]
  //: joint g20 (w28) @(254, 129) /w:[ 1 2 -1 4 ]
  mux g32 (.I0(w19), .I1(w5), .S(Cin), .Z(w31));   //: @(175,357) /sn:0 /delay:" 3 3" /w:[ 1 0 11 0 ] /ss:0 /do:0
  FA g0 (.A(w8), .B(w3), .Cin(w4), .Cout(w7), .S(w0));   //: @(438, 142) /sz:(61, 47) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Lo0<1 Bo0<1 ]
  tran g15(.Z(w23), .I(A[1]));   //: @(343,53) /sn:0 /R:1 /w:[ 3 4 3 ] /ss:1
  //: output g38 (S) @(318,495) /sn:0 /w:[ 1 ]
  mux g27 (.I0(w0), .I1(w1), .S(Cin), .Z(w6));   //: @(460,349) /sn:0 /delay:" 3 3" /w:[ 0 0 0 0 ] /ss:0 /do:0
  concat g37 (.I0(w6), .I1(w11), .I2(w29), .I3(w31), .Z(S));   //: @(310,446) /sn:0 /R:3 /w:[ 1 1 1 1 0 ] /dr:0
  tran g13(.Z(w32), .I(B[3]));   //: @(176,84) /sn:0 /R:1 /w:[ 3 8 7 ] /ss:1

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 {0}(116,382)(116,478)(272,478)(272,425)(215,425)(215,363)(302,363)(302,310){1}
wire [3:0] w0;    //: /sn:0 {0}(326,117)(326,211)(330,211)(330,221){1}
wire w1;    //: /sn:0 {0}(431,215)(612,215)(612,286)(465,286)(465,261)(376,261){1}
wire w2;    //: /sn:0 {0}(158,242)(158,338)(195,338)(195,271)(235,271){1}
wire [3:0] w5;    //: /sn:0 {0}(220,100)(220,211)(277,211)(277,221){1}
//: enddecls

  led g4 (.I(w2));   //: @(158,235) /sn:0 /w:[ 0 ] /type:0
  //: switch g3 (w1) @(414,215) /sn:0 /w:[ 0 ] /st:1
  //: dip g2 (w0) @(326,107) /sn:0 /w:[ 0 ] /st:5
  //: dip g1 (w5) @(220,90) /sn:0 /w:[ 0 ] /st:10
  led g5 (.I(w4));   //: @(116,375) /sn:0 /w:[ 0 ] /type:3
  CSA g0 (.B(w0), .A(w5), .Cin(w1), .Cout(w2), .S(w4));   //: @(236, 222) /sz:(139, 87) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule
