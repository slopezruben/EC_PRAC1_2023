//: version "1.8.7"

module CPA16(Cout, A, B, Cin, S);
//: interface  /sz:(149, 111) /bd:[ Ti0>A[15:0](44/149) Ti1>B[15:0](113/149) Ri0>Cin(42/111) Lo0<Cout(52/111) Bo0<S[15:0](69/149) ]
input [15:0] B;    //: /sn:0 {0}(-33,68)(129,68){1}
//: {2}(130,68)(300,68){3}
//: {4}(301,68)(479,68){5}
//: {6}(480,68)(668,68){7}
//: {8}(669,68)(694,68){9}
input [15:0] A;    //: /sn:0 {0}(36,31)(86,31){1}
//: {2}(87,31)(256,31){3}
//: {4}(257,31)(434,31){5}
//: {6}(435,31)(625,31){7}
//: {8}(626,31)(689,31){9}
input Cin;    //: /sn:0 {0}(796,173)(726,173)(726,171)(716,171){1}
output Cout;    //: /sn:0 {0}(26,315)(12,315)(12,191)(33,191){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(703,304)(883,304)(883,357)(846,357)(846,372)(856,372){1}
wire [3:0] w6;    //: /sn:0 {0}(435,149)(435,35){1}
wire w13;    //: /sn:0 {0}(204,184)(186,184)(186,183)(176,183){1}
wire [3:0] w16;    //: /sn:0 {0}(86,156)(86,43)(87,43)(87,35){1}
wire w7;    //: /sn:0 {0}(525,176)(563,176)(563,179)(573,179){1}
wire [3:0] w4;    //: /sn:0 {0}(609,224)(609,319)(697,319){1}
wire [3:0] w0;    //: /sn:0 {0}(670,144)(670,80)(669,80)(669,72){1}
wire [3:0] w19;    //: /sn:0 {0}(64,236)(64,289)(697,289){1}
wire [3:0] w10;    //: /sn:0 {0}(301,149)(301,72){1}
wire [3:0] w1;    //: /sn:0 {0}(626,144)(626,35){1}
wire w8;    //: /sn:0 {0}(382,184)(357,184)(357,176)(347,176){1}
wire [3:0] w14;    //: /sn:0 {0}(235,229)(235,299)(697,299){1}
wire [3:0] w11;    //: /sn:0 {0}(257,149)(257,35){1}
wire [3:0] w15;    //: /sn:0 {0}(130,156)(130,72){1}
wire [3:0] w5;    //: /sn:0 {0}(479,149)(479,78)(480,78)(480,72){1}
wire [3:0] w9;    //: /sn:0 {0}(413,229)(413,309)(697,309){1}
//: enddecls

  tran g8(.Z(w0), .I(B[3:0]));   //: @(669,66) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  //: output g4 (Cout) @(23,315) /sn:0 /w:[ 0 ]
  CPA4 g3 (.A(w16), .B(w15), .Cin(w13), .Cout(Cout), .S(w19));   //: @(34, 157) /sz:(141, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  concat g16 (.I0(w4), .I1(w9), .I2(w14), .I3(w19), .Z(S));   //: @(702,304) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  tran g17(.Z(w1), .I(A[3:0]));   //: @(626,29) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  CPA4 g2 (.A(w11), .B(w10), .Cin(w8), .Cout(w13), .S(w14));   //: @(205, 150) /sz:(141, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  CPA4 g1 (.A(w6), .B(w5), .Cin(w7), .Cout(w8), .S(w9));   //: @(383, 150) /sz:(141, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<0 Bo0<0 ]
  tran g10(.Z(w5), .I(B[7:4]));   //: @(480,66) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g6 (A) @(34,31) /sn:0 /w:[ 0 ]
  //: input g7 (B) @(-35,68) /sn:0 /w:[ 0 ]
  tran g9(.Z(w6), .I(A[7:4]));   //: @(435,29) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g12(.Z(w10), .I(B[11:8]));   //: @(301,66) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g14(.Z(w15), .I(B[15:12]));   //: @(130,66) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g5 (Cin) @(798,173) /sn:0 /R:2 /w:[ 0 ]
  tran g11(.Z(w11), .I(A[11:8]));   //: @(257,29) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  CPA4 g0 (.A(w1), .B(w0), .Cin(Cin), .Cout(w7), .S(w4));   //: @(574, 145) /sz:(141, 78) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  //: output g15 (S) @(853,372) /sn:0 /w:[ 1 ]
  tran g13(.Z(w16), .I(A[15:12]));   //: @(87,29) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule

module HA(S, B, C, A);
//: interface  /sz:(40, 40) /bd:[ Ti0>B(28/40) Ti1>A(8/40) Lo0<C(30/40) Bo0<S(17/40) ]
input B;    //: /sn:0 /dp:1 {0}(305,29)(207,29)(207,97){1}
//: {2}(209,99)(222,99)(222,93)(324,93){3}
//: {4}(207,101)(207,116)(197,116){5}
input A;    //: /sn:0 /dp:1 {0}(134,52)(171,52){1}
//: {2}(175,52)(195,52)(195,61)(231,61)(231,24)(305,24){3}
//: {4}(173,54)(173,71)(245,71){5}
output C;    //: /sn:0 /dp:1 {0}(345,91)(377,91){1}
output S;    //: /sn:0 /dp:1 {0}(326,27)(351,27){1}
wire w2;    //: /sn:0 {0}(261,71)(298,71)(298,88)(324,88){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(316,27) /sn:0 /delay:" 5" /w:[ 3 0 0 ]
  //: joint g8 (A) @(173, 52) /w:[ 2 -1 1 4 ]
  and g3 (.I0(w2), .I1(B), .Z(C));   //: @(335,91) /sn:0 /delay:" 4" /w:[ 1 3 0 ]
  //: output g2 (S) @(348,27) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(195,116) /sn:0 /w:[ 5 ]
  //: joint g6 (B) @(207, 99) /w:[ 2 1 -1 4 ]
  not g7 (.I(A), .Z(w2));   //: @(251,71) /sn:0 /w:[ 5 0 ]
  //: output g5 (C) @(374,91) /sn:0 /w:[ 1 ]
  //: input g0 (A) @(132,52) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire w7;    //: /sn:0 {0}(479,232)(479,217)(410,217){1}
wire [15:0] w4;    //: /sn:0 {0}(373,70)(373,174){1}
wire w0;    //: /sn:0 {0}(184,228)(184,238)(199,238)(199,227)(259,227){1}
wire [15:0] w1;    //: /sn:0 {0}(143,363)(143,373)(158,373)(158,385)(222,385)(222,308)(329,308)(329,287){1}
wire [15:0] w5;    //: /sn:0 {0}(241,89)(241,164)(304,164)(304,174){1}
//: enddecls

  led g4 (.I(w0));   //: @(184,221) /sn:0 /w:[ 0 ] /type:0
  //: switch g3 (w7) @(479,246) /sn:0 /R:1 /w:[ 0 ] /st:0
  //: dip g2 (w4) @(373,60) /sn:0 /w:[ 0 ] /st:3
  //: dip g1 (w5) @(241,79) /sn:0 /w:[ 0 ] /st:4
  led g5 (.I(w1));   //: @(143,356) /sn:0 /w:[ 0 ] /type:2
  CPA16 g0 (.A(w5), .B(w4), .Cin(w7), .Cout(w0), .S(w1));   //: @(260, 175) /sz:(149, 111) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule
