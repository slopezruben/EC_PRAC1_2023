//: version "1.8.7"

module RCA_2bits(M, B, A);
//: interface  /sz:(72, 50) /bd:[ Ti0>A[1:0](14/72) Ti1>B[1:0](41/72) Bo0<M[3:0](24/72) ]
output [3:0] M;    //: /sn:0 {0}(229,415)(229,343)(95,343)(95,325){1}
input [1:0] B;    //: /sn:0 {0}(366,89)(347,89){1}
//: {2}(346,89)(174,89){3}
//: {4}(173,89)(153,89)(153,83){5}
input [1:0] A;    //: /sn:0 {0}(328,53)(304,53){1}
//: {2}(303,53)(233,53){3}
//: {4}(232,53)(203,53)(203,66){5}
wire w7;    //: /sn:0 {0}(199,141)(199,157)(216,157)(216,167){1}
wire w0;    //: /sn:0 {0}(236,167)(236,140){1}
wire w3;    //: /sn:0 {0}(225,209)(225,292)(100,292)(100,319){1}
wire w12;    //: /sn:0 {0}(109,255)(109,279)(90,279)(90,319){1}
wire w10;    //: /sn:0 {0}(91,244)(80,244)(80,319){1}
wire w1;    //: /sn:0 {0}(110,319)(110,299)(346,299)(346,176){1}
wire w8;    //: /sn:0 {0}(304,57)(304,67)(319,67){1}
//: {2}(323,67)(343,67)(343,155){3}
//: {4}(321,69)(321,79)(201,79)(201,120){5}
wire w14;    //: /sn:0 {0}(91,180)(91,203)(100,203)(100,213){1}
wire w2;    //: /sn:0 {0}(207,198)(120,198)(120,213){1}
wire w11;    //: /sn:0 {0}(233,57)(233,64){1}
//: {2}(231,66)(88,66)(88,159){3}
//: {4}(233,68)(233,119){5}
wire w5;    //: /sn:0 {0}(174,93)(174,101)(176,101){1}
//: {2}(180,101)(196,101)(196,120){3}
//: {4}(178,103)(178,113)(93,113)(93,159){5}
wire w9;    //: /sn:0 {0}(347,93)(347,101)(348,101)(348,127){1}
//: {2}(346,129)(340,129)(340,115)(238,115)(238,119){3}
//: {4}(348,131)(348,155){5}
//: enddecls

  and g4 (.I0(w8), .I1(w9), .Z(w1));   //: @(346,166) /sn:0 /R:3 /delay:" 4" /w:[ 3 5 1 ]
  //: joint g8 (w9) @(348, 129) /w:[ -1 1 2 4 ]
  tran g3(.Z(w11), .I(A[1]));   //: @(233,51) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  concat g16 (.I0(w1), .I1(w3), .I2(w12), .I3(w10), .Z(M));   //: @(95,324) /sn:0 /R:3 /w:[ 0 1 1 1 1 ] /dr:1
  //: output g17 (M) @(229,412) /sn:0 /R:3 /w:[ 0 ]
  //: input g2 (B) @(368,89) /sn:0 /R:2 /w:[ 0 ]
  //: input g1 (A) @(330,53) /sn:0 /R:2 /w:[ 0 ]
  //: comment g18 /dolink:0 /link:"" @(364,169) /sn:0 /R:3
  //: /line:"a0 * b0"
  //: /end
  //: joint g10 (w8) @(321, 67) /w:[ 2 -1 1 4 ]
  tran g6(.Z(w9), .I(B[0]));   //: @(347,87) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  tran g7(.Z(w8), .I(A[0]));   //: @(304,51) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  and g9 (.I0(w5), .I1(w8), .Z(w7));   //: @(199,131) /sn:0 /R:3 /delay:" 4" /w:[ 3 5 0 ]
  HA g12 (.A(w14), .B(w2), .C(w10), .S(w12));   //: @(92, 214) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  and g5 (.I0(w11), .I1(w9), .Z(w0));   //: @(236,130) /sn:0 /R:3 /delay:" 4" /w:[ 5 3 1 ]
  tran g11(.Z(w5), .I(B[1]));   //: @(174,87) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  //: joint g14 (w5) @(178, 101) /w:[ 2 -1 1 4 ]
  //: comment g19 /dolink:0 /link:"" @(256,136) /sn:0 /R:3
  //: /line:"a1 * b0"
  //: /end
  //: comment g21 /dolink:0 /link:"" @(36,186) /sn:0 /R:3
  //: /line:"a1 * b1"
  //: /end
  //: comment g20 /dolink:0 /link:"" @(157,161) /sn:0 /R:3
  //: /line:"a0 * b1"
  //: /end
  HA g0 (.A(w7), .B(w0), .C(w2), .S(w3));   //: @(208, 168) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Lo0<0 Bo0<0 ]
  //: joint g15 (w11) @(233, 66) /w:[ -1 1 2 4 ]
  and g13 (.I0(w11), .I1(w5), .Z(w14));   //: @(91,170) /sn:0 /R:3 /delay:" 4" /w:[ 3 5 0 ]

endmodule

module main;    //: root_module
wire [1:0] w3;    //: /sn:0 {0}(329,62)(329,139)(298,139)(298,149){1}
wire [3:0] w1;    //: /sn:0 {0}(453,217)(453,277)(323,277)(323,223)(281,223)(281,201){1}
wire [1:0] w2;    //: /sn:0 {0}(235,60)(235,139)(271,139)(271,149){1}
//: enddecls

  led g3 (.I(w1));   //: @(453,210) /sn:0 /w:[ 0 ] /type:3
  //: dip g2 (w3) @(329,52) /sn:0 /w:[ 0 ] /st:3
  //: dip g1 (w2) @(235,50) /sn:0 /w:[ 0 ] /st:3
  RCA_2bits g0 (.B(w3), .A(w2), .M(w1));   //: @(257, 150) /sz:(72, 50) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]

endmodule
