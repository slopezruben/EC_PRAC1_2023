//: version "1.8.7"

module HA(S, B, C, A);
//: interface  /sz:(40, 40) /bd:[ Ti0>A(8/40) Ti1>B(28/40) Lo0<C(30/40) Bo0<S(17/40) ]
input B;    //: /sn:0 {0}(305,29)(207,29)(207,97){1}
//: {2}(209,99)(222,99)(222,93)(324,93){3}
//: {4}(207,101)(207,116)(197,116){5}
input A;    //: /sn:0 /dp:1 {0}(305,24)(225,24)(225,61)(189,61)(189,51){1}
//: {2}(191,49)(199,49)(199,88)(324,88){3}
//: {4}(189,47)(189,40)(177,40){5}
output C;    //: /sn:0 /dp:1 {0}(345,91)(377,91){1}
output S;    //: /sn:0 /dp:1 {0}(326,27)(351,27){1}
//: enddecls

  xor g4 (.I0(A), .I1(B), .Z(S));   //: @(316,27) /sn:0 /delay:" 5" /w:[ 0 0 0 ]
  and g3 (.I0(A), .I1(B), .Z(C));   //: @(335,91) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: output g2 (S) @(348,27) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(195,116) /sn:0 /w:[ 5 ]
  //: joint g6 (B) @(207, 99) /w:[ 2 1 -1 4 ]
  //: joint g7 (A) @(189, 49) /w:[ 2 4 -1 1 ]
  //: output g5 (C) @(374,91) /sn:0 /w:[ 1 ]
  //: input g0 (A) @(175,40) /sn:0 /w:[ 5 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(362,128)(362,113)(338,113)(338,103){1}
wire w7;    //: /sn:0 {0}(225,161)(310,161)(310,92)(320,92){1}
wire w4;    //: /sn:0 {0}(267,45)(267,51)(329,51)(329,61){1}
wire w5;    //: /sn:0 {0}(411,37)(411,51)(349,51)(349,61){1}
//: enddecls

  led g4 (.I(w7));   //: @(218,161) /sn:0 /R:1 /w:[ 0 ] /type:0
  led g3 (.I(w6));   //: @(362,135) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: switch g2 (w5) @(411,24) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: switch g1 (w4) @(267,32) /sn:0 /R:3 /w:[ 0 ] /st:0
  HA g0 (.B(w5), .A(w4), .C(w7), .S(w6));   //: @(321, 62) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]

endmodule
