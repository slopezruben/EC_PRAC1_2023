//: version "1.8.7"

module CPA4_alt(A, Cout, Cin, B, S);
//: interface  /sz:(141, 78) /bd:[ Ti0>B[3:0](96/141) Ti1>A[3:0](52/141) Ri0>Cin(26/78) Lo0<Cout(34/78) Bo0<S[3:0](30/141) ]
input [3:0] B;    //: /sn:0 {0}(96,106)(215,106){1}
//: {2}(216,106)(353,106){3}
//: {4}(354,106)(487,106){5}
//: {6}(488,106)(620,106){7}
//: {8}(621,106)(753,106){9}
input [3:0] A;    //: /sn:0 {0}(96,41)(191,41){1}
//: {2}(192,41)(328,41){3}
//: {4}(329,41)(463,41){5}
//: {6}(464,41)(596,41){7}
//: {8}(597,41)(745,41){9}
input Cin;    //: /sn:0 {0}(752,140)(776,140)(776,254)(655,254)(655,244){1}
output Cout;    //: /sn:0 /dp:1 {0}(283,218)(306,218)(306,203)(188,203)(188,187)(110,187)(110,421)(89,421){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(713,352)(762,352)(762,433)(772,433){1}
wire w13;    //: /sn:0 {0}(423,194)(444,194)(444,347)(707,347){1}
wire w6;    //: /sn:0 {0}(524,181)(464,181)(464,45){1}
wire w7;    //: /sn:0 {0}(635,215)(597,215)(597,45){1}
wire w4;    //: /sn:0 {0}(241,233)(192,233)(192,45){1}
wire w0;    //: /sn:0 {0}(381,184)(354,184)(354,110){1}
wire w3;    //: /sn:0 {0}(381,198)(329,198)(329,45){1}
wire w18;    //: /sn:0 {0}(566,186)(580,186)(580,242)(412,242)(412,223)(397,223)(397,213){1}
wire w12;    //: /sn:0 {0}(677,225)(694,225)(694,367)(707,367){1}
wire w19;    //: /sn:0 {0}(677,234)(687,234)(687,272)(540,272)(540,196){1}
wire w10;    //: /sn:0 {0}(635,229)(621,229)(621,110){1}
wire w1;    //: /sn:0 /dp:1 {0}(216,110)(216,219)(241,219){1}
wire w17;    //: /sn:0 {0}(566,177)(587,177)(587,357)(707,357){1}
wire w14;    //: /sn:0 {0}(423,203)(433,203)(433,274)(272,274)(272,258)(257,258)(257,248){1}
wire w5;    //: /sn:0 {0}(524,167)(488,167)(488,110){1}
wire w9;    //: /sn:0 {0}(283,229)(314,229)(314,337)(707,337){1}
//: enddecls

  //: input g4 (A) @(747,41) /sn:0 /R:2 /w:[ 9 ]
  tran g8(.Z(w5), .I(B[1]));   //: @(488,104) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: output g16 (Cout) @(92,421) /sn:0 /R:2 /w:[ 1 ]
  FA_alt g3 (.B(w10), .A(w7), .Ci(Cin), .Co(w19), .S(w12));   //: @(636, 203) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Bi0>1 Ro0<0 Ro1<0 ]
  //: input g17 (Cin) @(750,140) /sn:0 /w:[ 0 ]
  FA_alt g2 (.B(w6), .A(w5), .Ci(w19), .Co(w18), .S(w17));   //: @(525, 155) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Bi0>1 Ro0<0 Ro1<0 ]
  FA_alt g1 (.B(w3), .A(w0), .Ci(w18), .Co(w14), .S(w13));   //: @(382, 172) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>0 Bi0>1 Ro0<0 Ro1<0 ]
  //: comment g18 /dolink:0 /link:"" @(24,-51) /sn:0
  //: /line:"import Tarea03.v"
  //: /end
  tran g10(.Z(w0), .I(B[2]));   //: @(354,104) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g6(.Z(w10), .I(B[0]));   //: @(621,104) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g7(.Z(w7), .I(A[0]));   //: @(597,39) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g9(.Z(w6), .I(A[1]));   //: @(464,39) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g12(.Z(w1), .I(B[3]));   //: @(216,104) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: input g5 (B) @(755,106) /sn:0 /R:2 /w:[ 9 ]
  tran g11(.Z(w3), .I(A[2]));   //: @(329,39) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: output g14 (S) @(769,433) /sn:0 /w:[ 1 ]
  concat g15 (.I0(w12), .I1(w17), .I2(w13), .I3(w9), .Z(S));   //: @(712,352) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  FA_alt g0 (.B(w4), .A(w1), .Ci(w14), .Co(Cout), .S(w9));   //: @(242, 207) /sz:(40, 40) /sn:0 /p:[ Li0>0 Li1>1 Bi0>1 Ro0<0 Ro1<0 ]
  tran g13(.Z(w4), .I(A[3]));   //: @(192,39) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule

module main;    //: root_module
wire [3:0] w6;    //: /sn:0 {0}(289,57)(289,124)(263,124)(263,134){1}
wire [3:0] w7;    //: /sn:0 {0}(154,348)(154,358)(169,358)(169,316)(229,316)(229,226)(197,226)(197,214){1}
wire w3;    //: /sn:0 {0}(166,169)(99,169)(99,134){1}
wire w0;    //: /sn:0 {0}(410,120)(420,120)(420,135)(319,135)(319,161)(309,161){1}
wire [3:0] w5;    //: /sn:0 {0}(146,42)(146,124)(219,124)(219,134){1}
//: enddecls

  led g4 (.I(w3));   //: @(99,127) /sn:0 /w:[ 1 ] /type:0
  //: switch g3 (w0) @(393,120) /sn:0 /w:[ 0 ] /st:1
  //: dip g2 (w6) @(289,47) /sn:0 /w:[ 0 ] /st:15
  //: dip g1 (w5) @(146,32) /sn:0 /w:[ 0 ] /st:15
  led g5 (.I(w7));   //: @(154,341) /sn:0 /w:[ 0 ] /type:2
  CPA4_alt g0 (.B(w6), .A(w5), .Cin(w0), .Cout(w3), .S(w7));   //: @(167, 135) /sz:(141, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]

endmodule
