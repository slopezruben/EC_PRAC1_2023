//: version "1.8.7"

module Logic4(g3, g1, p1, g0, p0, C2, g2, p3, C1, C4, p2, C3, GG, Cin, PG);
//: interface  /sz:(514, 61) /bd:[ Ti0>p3(25/514) Ti1>g3(52/514) Ti2>p2(157/514) Ti3>g2(185/514) Ti4>p1(284/514) Ti5>g1(318/514) Ti6>p0(419/514) Ti7>g0(462/514) Ri0>Cin(28/61) To0<C3(121/514) To1<C2(251/514) To2<C1(387/514) Lo0<C4(28/61) Bo0<PG(69/514) Bo1<GG(48/514) ]
input g3;    //: /sn:0 {0}(73,363)(206,363)(206,283){1}
//: {2}(208,281)(228,281){3}
//: {4}(232,281)(454,281)(454,291)(514,291){5}
//: {6}(230,283)(230,406)(335,406){7}
//: {8}(204,281)(194,281)(194,282)(187,282){9}
input g2;    //: /sn:0 {0}(143,342)(214,342)(214,191){1}
//: {2}(216,189)(231,189){3}
//: {4}(235,189)(266,189){5}
//: {6}(270,189)(458,189){7}
//: {8}(268,191)(268,396)(335,396){9}
//: {10}(233,191)(233,438)(261,438){11}
//: {12}(212,189)(198,189)(198,191)(194,191){13}
output GG;    //: /sn:0 {0}(23,333)(33,333)(33,348)(16,348)(16,356)(52,356){1}
input g1;    //: /sn:0 {0}(130,288)(225,288)(225,137){1}
//: {2}(227,135)(245,135){3}
//: {4}(247,133)(247,127)(468,127){5}
//: {6}(247,137)(247,202)(284,202){7}
//: {8}(223,135)(212,135)(212,129)(200,129){9}
//: {10}(196,129)(184,129){11}
//: {12}(198,131)(198,401)(335,401){13}
output C3;    //: /sn:0 /dp:1 {0}(479,196)(520,196)(520,189)(531,189){1}
output PG;    //: /sn:0 /dp:1 {0}(83,166)(71,166)(71,125)(51,125){1}
input p3;    //: /sn:0 {0}(399,245)(176,245)(176,244)(166,244){1}
//: {2}(164,242)(164,68)(117,68){3}
//: {4}(164,246)(164,315){5}
//: {6}(166,317)(187,317){7}
//: {8}(191,317)(214,317){9}
//: {10}(218,317)(315,317){11}
//: {12}(319,317)(340,317){13}
//: {14}(344,317)(392,317){15}
//: {16}(342,319)(342,418)(251,418)(251,433)(261,433){17}
//: {18}(317,319)(317,363)(324,363){19}
//: {20}(328,363)(349,363){21}
//: {22}(326,361)(326,173)(104,173){23}
//: {24}(216,319)(216,347)(143,347){25}
//: {26}(189,315)(189,298)(130,298){27}
//: {28}(162,317)(149,317){29}
output C4;    //: /sn:0 /dp:1 {0}(535,301)(582,301)(582,294)(585,294){1}
output C2;    //: /sn:0 /dp:1 {0}(489,132)(540,132)(540,142)(547,142){1}
input Cin;    //: /sn:0 /dp:1 {0}(392,297)(364,297)(364,45){1}
//: {2}(366,43)(385,43)(385,25)(430,25){3}
//: {4}(362,43)(348,43){5}
//: {6}(344,43)(298,43){7}
//: {8}(294,43)(232,43)(232,44)(194,44){9}
//: {10}(296,45)(296,116)(346,116){11}
//: {12}(346,45)(346,148)(372,148)(372,235)(399,235){13}
input p2;    //: /sn:0 {0}(117,63)(209,63)(209,205){1}
//: {2}(211,207)(232,207){3}
//: {4}(236,207)(284,207){5}
//: {6}(234,209)(234,228)(244,228){7}
//: {8}(248,228)(261,228){9}
//: {10}(265,228)(279,228){11}
//: {12}(283,228)(303,228){13}
//: {14}(307,228)(350,228){15}
//: {16}(305,230)(305,358)(349,358){17}
//: {18}(281,230)(281,250)(399,250){19}
//: {20}(263,230)(263,255){21}
//: {22}(261,257)(251,257)(251,293)(130,293){23}
//: {24}(263,259)(263,312)(392,312){25}
//: {26}(246,226)(246,168)(104,168){27}
//: {28}(207,207)(201,207)(201,209)(195,209){29}
input p1;    //: /sn:0 {0}(117,58)(214,58)(214,150){1}
//: {2}(216,152)(227,152)(227,158)(236,158){3}
//: {4}(240,158)(251,158){5}
//: {6}(255,158)(271,158)(271,159)(288,159){7}
//: {8}(253,156)(253,121)(346,121){9}
//: {10}(253,160)(253,223)(350,223){11}
//: {12}(238,160)(238,172){13}
//: {14}(236,174)(227,174)(227,163)(104,163){15}
//: {16}(238,176)(238,307)(244,307){17}
//: {18}(248,307)(392,307){19}
//: {20}(246,309)(246,353)(349,353){21}
//: {22}(212,152)(193,152){23}
input p0;    //: /sn:0 {0}(104,158)(161,158)(161,110)(229,110)(229,96){1}
//: {2}(231,94)(279,94){3}
//: {4}(283,94)(304,94){5}
//: {6}(308,94)(387,94){7}
//: {8}(391,94)(424,94)(424,30)(430,30){9}
//: {10}(389,96)(389,240)(399,240){11}
//: {12}(306,96)(306,111)(346,111){13}
//: {14}(281,96)(281,302)(392,302){15}
//: {16}(227,94)(197,94)(197,95)(190,95){17}
input g0;    //: /sn:0 /dp:1 {0}(117,53)(236,53)(236,73){1}
//: {2}(238,75)(269,75){3}
//: {4}(273,75)(288,75){5}
//: {6}(292,75)(309,75){7}
//: {8}(313,75)(387,75)(387,49)(500,49){9}
//: {10}(311,77)(311,218)(350,218){11}
//: {12}(290,77)(290,348)(349,348){13}
//: {14}(271,77)(271,154)(288,154){15}
//: {16}(234,75)(216,75)(216,76)(190,76){17}
output C1;    //: /sn:0 {0}(564,35)(543,35)(543,47)(521,47){1}
wire w16;    //: /sn:0 {0}(73,358)(95,358)(95,344)(122,344){1}
wire w50;    //: /sn:0 {0}(413,307)(493,307)(493,296)(514,296){1}
wire w59;    //: /sn:0 {0}(282,436)(503,436)(503,306)(514,306){1}
wire w4;    //: /sn:0 {0}(73,348)(86,348)(86,61)(96,61){1}
wire w0;    //: /sn:0 {0}(73,353)(99,353)(99,293)(109,293){1}
wire w1;    //: /sn:0 {0}(514,311)(451,311)(451,381)(385,381)(385,401)(356,401){1}
wire w53;    //: /sn:0 {0}(370,355)(473,355)(473,345)(497,345)(497,301)(514,301){1}
wire w44;    //: /sn:0 {0}(371,223)(448,223)(448,204)(458,204){1}
wire w41;    //: /sn:0 {0}(305,205)(392,205)(392,194)(458,194){1}
wire w2;    //: /sn:0 {0}(451,28)(490,28)(490,44)(500,44){1}
wire w47;    //: /sn:0 {0}(420,242)(438,242)(438,199)(458,199){1}
wire w38;    //: /sn:0 {0}(367,116)(402,116)(402,132)(468,132){1}
wire w5;    //: /sn:0 {0}(309,157)(448,157)(448,137)(468,137){1}
//: enddecls

  //: joint g75 (p2) @(263, 257) /w:[ -1 21 22 24 ]
  //: joint g4 (g1) @(247, 135) /w:[ -1 4 3 6 ]
  //: joint g44 (p0) @(306, 94) /w:[ 6 -1 5 12 ]
  //: input g8 (g3) @(185,282) /sn:0 /w:[ 9 ]
  //: input g47 (g1) @(182,129) /sn:0 /w:[ 11 ]
  //: input g3 (p1) @(191,152) /sn:0 /w:[ 23 ]
  or g16 (.I0(w2), .I1(g0), .Z(C1));   //: @(511,47) /sn:0 /delay:" 4" /w:[ 1 9 1 ]
  and g26 (.I0(g0), .I1(p1), .Z(w5));   //: @(299,157) /sn:0 /delay:" 4" /w:[ 15 7 0 ]
  or g17 (.I0(g1), .I1(w38), .I2(w5), .Z(C2));   //: @(479,132) /sn:0 /delay:" 4" /w:[ 5 1 1 0 ]
  //: input g2 (g0) @(188,76) /sn:0 /w:[ 17 ]
  //: joint g74 (p3) @(189, 317) /w:[ 8 26 7 -1 ]
  and g30 (.I0(Cin), .I1(p0), .I2(p3), .I3(p2), .Z(w47));   //: @(410,242) /sn:0 /delay:" 4" /w:[ 13 11 0 19 0 ]
  //: joint g77 (g0) @(236, 75) /w:[ 2 1 16 -1 ]
  //: input g1 (p0) @(188,95) /sn:0 /w:[ 17 ]
  //: joint g60 (p2) @(305, 228) /w:[ 14 -1 13 16 ]
  and g29 (.I0(g0), .I1(p1), .I2(p2), .Z(w44));   //: @(361,223) /sn:0 /delay:" 4" /w:[ 11 11 15 0 ]
  //: joint g51 (p0) @(389, 94) /w:[ 8 -1 7 10 ]
  or g18 (.I0(g2), .I1(w41), .I2(w47), .I3(w44), .Z(C3));   //: @(469,196) /sn:0 /delay:" 4" /w:[ 7 1 1 1 0 ]
  //: joint g70 (p3) @(326, 363) /w:[ 20 22 19 -1 ]
  //: joint g65 (p3) @(342, 317) /w:[ 14 -1 13 16 ]
  //: output g10 (C2) @(544,142) /sn:0 /w:[ 1 ]
  //: joint g64 (g3) @(230, 281) /w:[ 4 -1 3 6 ]
  //: joint g49 (p2) @(234, 207) /w:[ 4 -1 3 6 ]
  //: joint g72 (p3) @(216, 317) /w:[ 10 -1 9 24 ]
  //: joint g50 (Cin) @(346, 43) /w:[ 5 -1 6 12 ]
  //: input g6 (g2) @(192,191) /sn:0 /w:[ 13 ]
  //: joint g58 (g0) @(290, 75) /w:[ 6 -1 5 12 ]
  //: joint g56 (p1) @(238, 158) /w:[ 4 -1 3 12 ]
  and g35 (.I0(p3), .I1(p2), .I2(p1), .I3(p0), .Z(PG));   //: @(93,166) /sn:0 /R:2 /delay:" 4" /w:[ 23 27 15 0 0 ]
  //: input g7 (p3) @(147,317) /sn:0 /w:[ 29 ]
  //: output g9 (C1) @(561,35) /sn:0 /w:[ 0 ]
  //: joint g68 (p1) @(238, 174) /w:[ -1 13 14 16 ]
  //: joint g73 (g2) @(214, 189) /w:[ 2 -1 12 1 ]
  //: joint g59 (p1) @(246, 307) /w:[ 18 -1 17 20 ]
  and g31 (.I0(Cin), .I1(p0), .I2(p1), .I3(p2), .I4(p3), .Z(w50));   //: @(403,307) /sn:0 /delay:" 4" /w:[ 0 15 19 25 15 0 ]
  //: joint g71 (g3) @(206, 281) /w:[ 2 -1 8 1 ]
  //: joint g67 (p0) @(229, 94) /w:[ 2 -1 16 1 ]
  //: joint g54 (Cin) @(364, 43) /w:[ 2 -1 4 1 ]
  //: joint g45 (Cin) @(296, 43) /w:[ 7 -1 8 10 ]
  and g36 (.I0(p3), .I1(g2), .Z(w16));   //: @(132,344) /sn:0 /R:2 /delay:" 4" /w:[ 25 0 1 ]
  and g33 (.I0(g2), .I1(g1), .I2(g3), .Z(w1));   //: @(346,401) /sn:0 /delay:" 4" /w:[ 9 13 7 1 ]
  //: joint g69 (p2) @(246, 228) /w:[ 8 26 7 -1 ]
  //: joint g66 (g2) @(233, 189) /w:[ 4 -1 3 10 ]
  //: output g12 (C4) @(582,294) /sn:0 /w:[ 1 ]
  //: joint g57 (p2) @(263, 228) /w:[ 10 -1 9 20 ]
  //: joint g46 (p1) @(253, 158) /w:[ 6 8 5 10 ]
  and g34 (.I0(p3), .I1(g2), .Z(w59));   //: @(272,436) /sn:0 /delay:" 4" /w:[ 17 11 0 ]
  and g28 (.I0(g1), .I1(p2), .Z(w41));   //: @(295,205) /sn:0 /delay:" 4" /w:[ 7 5 0 ]
  //: input g5 (p2) @(193,209) /sn:0 /w:[ 29 ]
  //: output g11 (C3) @(528,189) /sn:0 /w:[ 1 ]
  //: output g14 (GG) @(26,333) /sn:0 /R:2 /w:[ 0 ]
  //: joint g61 (p3) @(317, 317) /w:[ 12 -1 11 18 ]
  or g19 (.I0(g3), .I1(w50), .I2(w53), .I3(w59), .I4(w1), .Z(C4));   //: @(525,301) /sn:0 /delay:" 4" /w:[ 5 1 1 1 0 0 ]
  //: joint g21 (p3) @(164, 244) /w:[ 1 2 -1 4 ]
  //: joint g79 (p2) @(209, 207) /w:[ 2 1 28 -1 ]
  //: joint g78 (p1) @(214, 152) /w:[ 2 1 22 -1 ]
  and g32 (.I0(g0), .I1(p1), .I2(p2), .I3(p3), .Z(w53));   //: @(360,355) /sn:0 /delay:" 4" /w:[ 13 21 17 21 0 ]
  or g20 (.I0(g3), .I1(w16), .I2(w0), .I3(w4), .Z(GG));   //: @(62,356) /sn:0 /R:2 /delay:" 4" /w:[ 0 0 0 0 1 ]
  //: joint g63 (g2) @(268, 189) /w:[ 6 -1 5 8 ]
  //: joint g43 (g0) @(271, 75) /w:[ 4 -1 3 14 ]
  and g38 (.I0(p3), .I1(p2), .I2(p1), .I3(g0), .Z(w4));   //: @(106,61) /sn:0 /R:2 /delay:" 4" /w:[ 3 0 0 0 1 ]
  //: input g0 (Cin) @(192,44) /sn:0 /w:[ 9 ]
  and g15 (.I0(Cin), .I1(p0), .Z(w2));   //: @(441,28) /sn:0 /delay:" 4" /w:[ 3 9 0 ]
  //: joint g48 (g0) @(311, 75) /w:[ 8 -1 7 10 ]
  and g27 (.I0(p0), .I1(Cin), .I2(p1), .Z(w38));   //: @(357,116) /sn:0 /delay:" 4" /w:[ 13 11 9 0 ]
  //: joint g62 (g1) @(198, 129) /w:[ 9 -1 10 12 ]
  and g37 (.I0(p3), .I1(p2), .I2(g1), .Z(w0));   //: @(119,293) /sn:0 /R:2 /delay:" 4" /w:[ 27 23 0 1 ]
  //: joint g80 (p3) @(164, 317) /w:[ 6 5 28 -1 ]
  //: joint g55 (p0) @(281, 94) /w:[ 4 -1 3 14 ]
  //: joint g76 (g1) @(225, 135) /w:[ 2 -1 8 1 ]
  //: joint g53 (p2) @(281, 228) /w:[ 12 -1 11 18 ]
  //: output g13 (PG) @(54,125) /sn:0 /R:2 /w:[ 1 ]

endmodule

module CLA4(S, B, Cin, A, Cout, GG, PG);
//: interface  /sz:(108, 57) /bd:[ Ti0>A[3:0](19/108) Ti1>B[3:0](76/108) Ri0>Cin(27/57) Lo0<Cout(28/57) Bo0<S[3:0](45/108) Bo1<PG(75/108) Bo2<GG(96/108) ]
input [3:0] B;    //: /sn:0 /dp:5 {0}(611,57)(588,57){1}
//: {2}(587,57)(447,57){3}
//: {4}(446,57)(316,57){5}
//: {6}(315,57)(183,57){7}
//: {8}(182,57)(56,57){9}
output GG;    //: /sn:0 {0}(131,375)(131,311)(168,311)(168,301){1}
input [3:0] A;    //: /sn:0 {0}(57,16)(151,16){1}
//: {2}(152,16)(282,16){3}
//: {4}(283,16)(415,16){5}
//: {6}(416,16)(552,16){7}
//: {8}(553,16)(621,16){9}
output PG;    //: /sn:0 {0}(170,374)(170,344)(189,344)(189,301){1}
input Cin;    //: /sn:0 {0}(705,180)(685,180)(685,178)(644,178){1}
//: {2}(640,178)(637,178)(637,149)(629,149){3}
//: {4}(642,180)(642,267)(635,267){5}
output Cout;    //: /sn:0 {0}(55,266)(43,266)(43,253)(109,253)(109,267)(119,267){1}
output [3:0] S;    //: /sn:0 {0}(649,341)(673,341)(673,409)(680,409){1}
wire w6;    //: /sn:0 {0}(445,119)(445,69)(447,69)(447,61){1}
wire w13;    //: /sn:0 {0}(283,120)(283,20){1}
wire w16;    //: /sn:0 {0}(306,181)(306,217)(305,217)(305,238){1}
wire w7;    //: /sn:0 {0}(413,119)(413,28)(416,28)(416,20){1}
wire w25;    //: /sn:0 /dp:1 {0}(507,238)(507,148)(485,148){1}
wire w0;    //: /sn:0 {0}(589,120)(589,69)(588,69)(588,61){1}
wire w3;    //: /sn:0 {0}(548,181)(548,228)(539,228)(539,238){1}
wire w22;    //: /sn:0 {0}(174,181)(174,210)(172,210)(172,238){1}
wire w20;    //: /sn:0 /dp:1 {0}(404,238)(404,180){1}
wire w12;    //: /sn:0 {0}(315,120)(315,69)(316,69)(316,61){1}
wire w18;    //: /sn:0 {0}(183,120)(183,61){1}
wire w19;    //: /sn:0 {0}(151,120)(151,28)(152,28)(152,20){1}
wire w10;    //: /sn:0 {0}(436,180)(436,228)(438,228)(438,238){1}
wire w23;    //: /sn:0 {0}(205,181)(205,326)(643,326){1}
wire w21;    //: /sn:0 {0}(142,181)(142,228)(145,228)(145,238){1}
wire w1;    //: /sn:0 {0}(557,120)(557,28)(553,28)(553,20){1}
wire w17;    //: /sn:0 {0}(337,181)(337,336)(643,336){1}
wire w27;    //: /sn:0 /dp:1 {0}(241,238)(241,149)(223,149){1}
wire w28;    //: /sn:0 /dp:1 {0}(277,238)(277,192)(274,192)(274,181){1}
wire w11;    //: /sn:0 {0}(467,180)(467,346)(643,346){1}
wire w2;    //: /sn:0 /dp:1 {0}(582,238)(582,192)(580,192)(580,181){1}
wire w5;    //: /sn:0 {0}(611,181)(611,356)(643,356){1}
wire w26;    //: /sn:0 /dp:1 {0}(371,238)(371,149)(355,149){1}
//: enddecls

  PFA g4 (.a(w19), .b(w18), .Ci(w27), .Si(w23), .Gi(w22), .Pi(w21));   //: @(122, 121) /sz:(100, 59) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<0 ]
  //: output g8 (S) @(677,409) /sn:0 /w:[ 1 ]
  PFA g3 (.a(w13), .b(w12), .Ci(w26), .Si(w17), .Gi(w16), .Pi(w28));   //: @(254, 121) /sz:(100, 59) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  tran g16(.Z(w13), .I(A[2]));   //: @(283,14) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g17(.Z(w18), .I(B[3]));   //: @(183,55) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  PFA g2 (.a(w7), .b(w6), .Ci(w25), .Si(w11), .Gi(w10), .Pi(w20));   //: @(384, 120) /sz:(100, 59) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Bo0<0 Bo1<0 Bo2<1 ]
  PFA g1 (.a(w1), .b(w0), .Ci(Cin), .Si(w5), .Gi(w2), .Pi(w3));   //: @(528, 121) /sz:(100, 59) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>3 Bo0<0 Bo1<1 Bo2<0 ]
  tran g18(.Z(w19), .I(A[3]));   //: @(152,14) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: input g10 (B) @(54,57) /sn:0 /w:[ 9 ]
  //: input g6 (Cin) @(707,180) /sn:0 /R:2 /w:[ 0 ]
  //: joint g7 (Cin) @(642, 178) /w:[ 1 -1 2 4 ]
  //: input g9 (A) @(55,16) /sn:0 /w:[ 0 ]
  tran g12(.Z(w1), .I(A[0]));   //: @(553,14) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  concat g5 (.I0(w5), .I1(w11), .I2(w17), .I3(w23), .Z(S));   //: @(648,341) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  tran g11(.Z(w0), .I(B[0]));   //: @(588,55) /sn:0 /R:1 /w:[ 1 2 1 ] /ss:1
  tran g14(.Z(w7), .I(A[1]));   //: @(416,14) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: output g19 (Cout) @(52,266) /sn:0 /w:[ 0 ]
  //: output g21 (GG) @(131,372) /sn:0 /R:3 /w:[ 0 ]
  //: output g20 (PG) @(170,371) /sn:0 /R:3 /w:[ 0 ]
  Logic4 g0 (.p3(w21), .g3(w22), .p2(w28), .g2(w16), .p1(w20), .g1(w10), .p0(w3), .g0(w2), .Cin(Cin), .C3(w27), .C2(w26), .C1(w25), .C4(Cout), .PG(PG), .GG(GG));   //: @(120, 239) /sz:(514, 61) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>0 Ti3>1 Ti4>0 Ti5>1 Ti6>1 Ti7>0 Ri0>5 To0<0 To1<0 To2<0 Lo0<1 Bo0<1 Bo1<1 ]
  tran g15(.Z(w12), .I(B[2]));   //: @(316,55) /sn:0 /R:1 /w:[ 1 6 5 ] /ss:1
  tran g13(.Z(w6), .I(B[1]));   //: @(447,55) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1

endmodule

module main;    //: root_module
wire [3:0] w7;    //: /sn:0 {0}(118,86)(118,191)(185,191)(185,201){1}
wire w4;    //: /sn:0 {0}(222,366)(222,313)(231,313)(231,288)(241,288)(241,260){1}
wire w0;    //: /sn:0 {0}(96,247)(96,257)(111,257)(111,230)(165,230){1}
wire w3;    //: /sn:0 /dp:1 {0}(275,229)(357,229)(357,258){1}
wire [3:0] w1;    //: /sn:0 /dp:1 {0}(242,201)(242,98)(310,98)(310,88){1}
wire w8;    //: /sn:0 {0}(270,309)(270,270)(262,270)(262,260){1}
wire [3:0] w5;    //: /sn:0 {0}(90,335)(90,345)(122,345)(122,275)(211,275)(211,260){1}
//: enddecls

  //: switch g4 (w3) @(357,272) /sn:0 /R:1 /w:[ 1 ] /st:0
  led g3 (.I(w0));   //: @(96,240) /sn:0 /w:[ 0 ] /type:0
  //: dip g2 (w1) @(310,78) /sn:0 /w:[ 1 ] /st:15
  //: dip g1 (w7) @(118,76) /sn:0 /w:[ 0 ] /st:1
  led g6 (.I(w8));   //: @(270,316) /sn:0 /R:2 /w:[ 0 ] /type:0
  led g7 (.I(w5));   //: @(90,328) /sn:0 /w:[ 0 ] /type:2
  led g5 (.I(w4));   //: @(222,373) /sn:0 /R:2 /w:[ 0 ] /type:0
  CLA4 g0 (.B(w1), .A(w7), .Cin(w3), .Cout(w0), .GG(w8), .PG(w4), .S(w5));   //: @(166, 202) /sz:(108, 57) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Bo0<1 Bo1<1 Bo2<1 ]

endmodule
