//: version "1.8.7"

module CSA16(A, Cout, Cin, S, B);
//: interface  /sz:(162, 100) /bd:[ Ti0>B[15:0](115/162) Ti1>A[15:0](34/162) Ri0>Cin(49/100) Lo0<Cout(46/100) Bo0<S[15:0](79/162) ]
input [15:0] B;    //: /sn:0 {0}(84,54)(244,54){1}
//: {2}(245,54)(414,54){3}
//: {4}(415,54)(587,54){5}
//: {6}(588,54)(789,54){7}
//: {8}(790,54)(825,54)(825,45){9}
input [15:0] A;    //: /sn:0 {0}(85,19)(189,19){1}
//: {2}(190,19)(361,19){3}
//: {4}(362,19)(537,19){5}
//: {6}(538,19)(738,19){7}
//: {8}(739,19)(813,19){9}
input Cin;    //: /sn:0 {0}(921,195)(848,195)(848,196)(838,196){1}
output Cout;    //: /sn:0 {0}(65,210)(140,210)(140,208)(150,208){1}
output [15:0] S;    //: /sn:0 {0}(851,242)(841,242)(841,257)(937,257)(937,286)(930,286)(930,305)(1014,305)(1014,399)(1006,399)(1006,389)(880,389){1}
wire [3:0] w6;    //: /sn:0 {0}(538,162)(538,23){1}
wire w13;    //: /sn:0 {0}(318,208)(301,208)(301,198)(291,198){1}
wire [3:0] w16;    //: /sn:0 {0}(192,158)(192,31)(190,31)(190,23){1}
wire [3:0] w4;    //: /sn:0 {0}(764,245)(764,404)(874,404){1}
wire [3:0] w0;    //: /sn:0 {0}(792,156)(792,66)(790,66)(790,58){1}
wire w3;    //: /sn:0 {0}(697,206)(647,206)(647,202)(637,202){1}
wire [3:0] w19;    //: /sn:0 {0}(217,247)(217,374)(874,374){1}
wire [3:0] w10;    //: /sn:0 {0}(413,158)(413,66)(415,66)(415,58){1}
wire [3:0] w1;    //: /sn:0 {0}(739,156)(739,23){1}
wire w8;    //: /sn:0 {0}(496,212)(469,212)(469,198)(459,198){1}
wire [3:0] w14;    //: /sn:0 {0}(385,247)(385,384)(874,384){1}
wire [3:0] w11;    //: /sn:0 {0}(360,158)(360,27)(362,27)(362,23){1}
wire [3:0] w15;    //: /sn:0 {0}(245,158)(245,58){1}
wire [3:0] w5;    //: /sn:0 {0}(591,162)(591,66)(588,66)(588,58){1}
wire [3:0] w9;    //: /sn:0 {0}(563,251)(563,394)(874,394){1}
//: enddecls

  //: input g4 (A) @(83,19) /sn:0 /w:[ 0 ]
  //: output g8 (Cout) @(68,210) /sn:0 /R:2 /w:[ 0 ]
  CSA g3 (.A(w16), .B(w15), .Cin(w13), .Cout(Cout), .S(w19));   //: @(151, 159) /sz:(139, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<0 ]
  tran g16(.Z(w1), .I(A[3:0]));   //: @(739,17) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g17(.Z(w0), .I(B[3:0]));   //: @(790,52) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  CSA g2 (.A(w11), .B(w10), .Cin(w8), .Cout(w13), .S(w14));   //: @(319, 159) /sz:(139, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  CSA g1 (.A(w6), .B(w5), .Cin(w3), .Cout(w8), .S(w9));   //: @(497, 163) /sz:(139, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  tran g10(.Z(w16), .I(A[15:12]));   //: @(190,17) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  concat g6 (.I0(w4), .I1(w9), .I2(w14), .I3(w19), .Z(S));   //: @(879,389) /sn:0 /w:[ 1 1 1 1 1 ] /dr:0
  //: input g7 (Cin) @(923,195) /sn:0 /R:2 /w:[ 0 ]
  //: output g9 (S) @(848,242) /sn:0 /w:[ 0 ]
  tran g12(.Z(w11), .I(A[11:8]));   //: @(362,17) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g5 (B) @(82,54) /sn:0 /w:[ 0 ]
  tran g11(.Z(w15), .I(B[15:12]));   //: @(245,52) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g14(.Z(w6), .I(A[7:4]));   //: @(538,17) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  CSA g0 (.A(w1), .B(w0), .Cin(Cin), .Cout(w3), .S(w4));   //: @(698, 157) /sz:(139, 87) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  tran g15(.Z(w5), .I(B[7:4]));   //: @(588,52) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g13(.Z(w10), .I(B[11:8]));   //: @(415,52) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 {0}(435,91)(435,168)(387,168)(387,178){1}
wire w4;    //: /sn:0 /dp:1 {0}(435,228)(507,228)(507,252){1}
wire [15:0] w3;    //: /sn:0 {0}(274,87)(274,168)(306,168)(306,178){1}
wire w2;    //: /sn:0 {0}(164,235)(164,243)(196,243)(196,225)(271,225){1}
wire [15:0] w5;    //: /sn:0 {0}(337,411)(337,421)(351,421)(351,280){1}
//: enddecls

  //: dip g4 (w3) @(274,77) /sn:0 /w:[ 0 ] /st:10
  led g3 (.I(w2));   //: @(164,228) /sn:0 /w:[ 0 ] /type:0
  //: switch g2 (w4) @(507,266) /sn:0 /R:1 /w:[ 1 ] /st:0
  led g1 (.I(w5));   //: @(337,404) /sn:0 /w:[ 0 ] /type:3
  //: dip g5 (w6) @(435,81) /sn:0 /w:[ 0 ] /st:170
  CSA16 g0 (.B(w6), .A(w3), .Cin(w4), .Cout(w2), .S(w5));   //: @(272, 179) /sz:(162, 100) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Lo0<1 Bo0<1 ]

endmodule
