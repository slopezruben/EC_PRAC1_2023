//: version "1.8.7"

module CPA4(A, Cout, Cin, S, B);
//: interface  /sz:(141, 78) /bd:[ Ti0>A[3:0](52/141) Ti1>B[3:0](96/141) Ri0>Cin(26/78) Lo0<Cout(34/78) Bo0<S[3:0](30/141) ]
input [3:0] B;    //: /sn:0 {0}(96,106)(215,106){1}
//: {2}(216,106)(353,106){3}
//: {4}(354,106)(487,106){5}
//: {6}(488,106)(620,106){7}
//: {8}(621,106)(753,106){9}
input [3:0] A;    //: /sn:0 {0}(96,41)(191,41){1}
//: {2}(192,41)(328,41){3}
//: {4}(329,41)(463,41){5}
//: {6}(464,41)(596,41){7}
//: {8}(597,41)(745,41){9}
input Cin;    //: /sn:0 {0}(752,140)(762,140)(762,155)(651,155)(651,164)(641,164){1}
output Cout;    //: /sn:0 /dp:1 {0}(177,209)(99,209)(99,421)(89,421){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(713,352)(762,352)(762,433)(772,433){1}
wire w16;    //: /sn:0 {0}(622,146)(622,118)(621,118)(621,110){1}
wire w13;    //: /sn:0 {0}(447,181)(382,181)(382,190)(372,190){1}
wire w6;    //: /sn:0 {0}(353,172)(353,118)(354,118)(354,110){1}
wire w7;    //: /sn:0 /dp:1 {0}(707,357)(473,357)(473,199){1}
wire w0;    //: /sn:0 {0}(194,185)(194,53)(192,53)(192,45){1}
wire w20;    //: /sn:0 {0}(707,347)(337,347)(337,214){1}
wire w18;    //: /sn:0 {0}(580,170)(518,170)(518,175)(508,175){1}
wire w10;    //: /sn:0 {0}(464,157)(464,45){1}
wire w21;    //: /sn:0 {0}(707,337)(203,337)(203,227){1}
wire w1;    //: /sn:0 {0}(219,185)(219,118)(216,118)(216,110){1}
wire w8;    //: /sn:0 {0}(311,196)(248,196)(248,203)(238,203){1}
wire w2;    //: /sn:0 /dp:1 {0}(707,367)(606,367)(606,188){1}
wire w11;    //: /sn:0 {0}(489,157)(489,118)(488,118)(488,110){1}
wire w15;    //: /sn:0 {0}(597,146)(597,45){1}
wire w5;    //: /sn:0 {0}(328,172)(328,53)(329,53)(329,45){1}
//: enddecls

  tran g8(.Z(w11), .I(B[1]));   //: @(488,104) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g4 (A) @(747,41) /sn:0 /R:2 /w:[ 9 ]
  //: output g16 (Cout) @(92,421) /sn:0 /R:2 /w:[ 1 ]
  FA g3 (.B(w16), .A(w15), .Cin(Cin), .Cout(w18), .S(w2));   //: @(581, 147) /sz:(59, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  //: input g17 (Cin) @(750,140) /sn:0 /w:[ 0 ]
  FA g2 (.B(w11), .A(w10), .Cin(w18), .Cout(w13), .S(w7));   //: @(448, 158) /sz:(59, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  FA g1 (.B(w6), .A(w5), .Cin(w13), .Cout(w8), .S(w20));   //: @(312, 173) /sz:(59, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  tran g10(.Z(w6), .I(B[2]));   //: @(354,104) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  tran g6(.Z(w16), .I(B[0]));   //: @(621,104) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g9(.Z(w10), .I(A[1]));   //: @(464,39) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g7(.Z(w15), .I(A[0]));   //: @(597,39) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g12(.Z(w1), .I(B[3]));   //: @(216,104) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g14 (S) @(769,433) /sn:0 /w:[ 1 ]
  tran g11(.Z(w5), .I(A[2]));   //: @(329,39) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: input g5 (B) @(755,106) /sn:0 /R:2 /w:[ 9 ]
  concat g15 (.I0(w2), .I1(w7), .I2(w20), .I3(w21), .Z(S));   //: @(712,352) /sn:0 /w:[ 0 0 0 0 0 ] /dr:0
  FA g0 (.B(w1), .A(w0), .Cin(w8), .Cout(Cout), .S(w21));   //: @(178, 186) /sz:(59, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 ]
  tran g13(.Z(w0), .I(A[3]));   //: @(192,39) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1

endmodule

module main;    //: root_module
wire [3:0] w6;    //: /sn:0 {0}(289,57)(289,124)(263,124)(263,134){1}
wire [3:0] w7;    //: /sn:0 {0}(154,348)(154,358)(169,358)(169,316)(229,316)(229,226)(197,226)(197,214){1}
wire w0;    //: /sn:0 {0}(410,120)(420,120)(420,135)(319,135)(319,161)(309,161){1}
wire w3;    //: /sn:0 {0}(166,169)(99,169)(99,134){1}
wire [3:0] w5;    //: /sn:0 {0}(146,42)(146,124)(219,124)(219,134){1}
//: enddecls

  led g4 (.I(w3));   //: @(99,127) /sn:0 /w:[ 1 ] /type:0
  //: switch g3 (w0) @(393,120) /sn:0 /w:[ 0 ] /st:1
  //: dip g2 (w6) @(289,47) /sn:0 /w:[ 0 ] /st:15
  //: dip g1 (w5) @(146,32) /sn:0 /w:[ 0 ] /st:15
  led g5 (.I(w7));   //: @(154,341) /sn:0 /w:[ 0 ] /type:2
  CPA4 g0 (.B(w6), .A(w5), .Cin(w0), .Cout(w3), .S(w7));   //: @(167, 135) /sz:(141, 78) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]

endmodule
