//: version "1.8.7"

module CLA16(S, PG, GG, Cin, A, Cout, B);
//: interface  /sz:(141, 84) /bd:[ Ti0>B[15:0](103/141) Ti1>A[15:0](31/141) Ri0>Cin(44/84) Lo0<Cout(39/84) Bo0<GG(125/141) Bo1<PG(104/141) Bo2<S[15:0](65/141) ]
input [15:0] B;    //: /sn:0 {0}(153,87)(265,87){1}
//: {2}(266,87)(415,87){3}
//: {4}(416,87)(489,87)(489,86)(610,86){5}
//: {6}(611,86)(766,86)(766,87)(776,87){7}
//: {8}(777,87)(806,87){9}
output GG;    //: /sn:0 {0}(259,429)(249,429)(249,414)(263,414)(263,380){1}
input [15:0] A;    //: /sn:0 {0}(152,43)(207,43){1}
//: {2}(208,43)(355,43){3}
//: {4}(356,43)(552,43){5}
//: {6}(553,43)(718,43){7}
//: {8}(719,43)(822,43){9}
output PG;    //: /sn:0 /dp:1 {0}(284,380)(284,431)(319,431){1}
input Cin;    //: /sn:0 {0}(730,346)(828,346)(828,208){1}
//: {2}(830,206)(898,206){3}
//: {4}(826,206)(818,206)(818,184)(810,184){5}
output Cout;    //: /sn:0 /dp:1 {0}(214,346)(186,346){1}
//: {2}(182,346)(175,346){3}
//: {4}(184,348)(184,358)(167,358)(167,345)(150,345){5}
output [15:0] S;    //: /sn:0 {0}(956,407)(878,407)(878,418)(868,418){1}
wire w13;    //: /sn:0 {0}(634,317)(634,261)(776,261)(776,215){1}
wire w16;    //: /sn:0 {0}(336,317)(336,274)(315,274)(315,187)(297,187){1}
wire w7;    //: /sn:0 /dp:1 {0}(372,317)(372,276)(415,276)(415,200){1}
wire w39;    //: /sn:0 {0}(187,188)(170,188)(170,168){1}
wire [3:0] w0;    //: /sn:0 {0}(720,156)(720,55)(719,55)(719,47){1}
wire [3:0] w22;    //: /sn:0 {0}(553,132)(553,47){1}
wire [3:0] w36;    //: /sn:0 {0}(207,159)(207,103)(208,103)(208,47){1}
wire [3:0] w3;    //: /sn:0 /dp:1 {0}(862,423)(579,423)(579,191){1}
wire [3:0] w29;    //: /sn:0 {0}(359,141)(359,55)(356,55)(356,47){1}
wire [3:0] w30;    //: /sn:0 {0}(416,141)(416,91){1}
wire [3:0] w37;    //: /sn:0 {0}(264,159)(264,99)(266,99)(266,91){1}
wire w42;    //: /sn:0 {0}(284,218)(284,307)(267,307)(267,317){1}
wire w12;    //: /sn:0 {0}(533,317)(533,251)(630,251)(630,191){1}
wire w18;    //: /sn:0 {0}(602,317)(602,293)(655,293)(655,160)(643,160){1}
wire [3:0] w23;    //: /sn:0 {0}(610,132)(610,98)(611,98)(611,90){1}
wire w10;    //: /sn:0 /dp:1 {0}(685,166)(685,185)(700,185){1}
wire [3:0] w1;    //: /sn:0 {0}(777,156)(777,91){1}
wire w32;    //: /sn:0 {0}(339,170)(318,170)(318,150){1}
wire [3:0] w8;    //: /sn:0 {0}(862,413)(385,413)(385,200){1}
wire w17;    //: /sn:0 {0}(466,317)(466,169)(449,169){1}
wire w14;    //: /sn:0 {0}(677,317)(677,278)(797,278)(797,215){1}
wire w11;    //: /sn:0 {0}(499,317)(499,228)(609,228)(609,191){1}
wire w41;    //: /sn:0 {0}(263,218)(263,307)(240,307)(240,317){1}
wire [3:0] w2;    //: /sn:0 /dp:1 {0}(862,433)(746,433)(746,215){1}
wire [3:0] w15;    //: /sn:0 {0}(862,403)(233,403)(233,218){1}
wire w5;    //: /sn:0 /dp:1 {0}(400,317)(400,292)(436,292)(436,200){1}
wire w9;    //: /sn:0 /dp:1 {0}(511,153)(511,161)(533,161){1}
//: enddecls

  CLA4 g4 (.B(w37), .A(w36), .Cin(w16), .Cout(w39), .GG(w42), .PG(w41), .S(w15));   //: @(188, 160) /sz:(108, 57) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<0 Bo1<0 Bo2<1 ]
  led g8 (.I(w10));   //: @(685,159) /sn:0 /w:[ 0 ] /type:0
  CLA4 g3 (.B(w30), .A(w29), .Cin(w17), .Cout(w32), .GG(w5), .PG(w7), .S(w8));   //: @(340, 142) /sz:(108, 57) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<0 Bo0<1 Bo1<1 Bo2<1 ]
  //: output g16 (S) @(953,407) /sn:0 /w:[ 0 ]
  tran g17(.Z(w36), .I(A[15:12]));   //: @(208,41) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  //: output g26 (PG) @(316,431) /sn:0 /w:[ 1 ]
  CLA4 g2 (.B(w23), .A(w22), .Cin(w18), .Cout(w9), .GG(w12), .PG(w11), .S(w3));   //: @(534, 133) /sz:(108, 57) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Bo2<1 ]
  tran g23(.Z(w30), .I(B[11:8]));   //: @(416,85) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  Logic4 g1 (.g0(w14), .p0(w13), .g1(w12), .p1(w11), .g2(w5), .p2(w7), .g3(w42), .p3(w41), .Cin(Cin), .C1(w18), .C2(w17), .C3(w16), .C4(Cout), .GG(GG), .PG(PG));   //: @(215, 318) /sz:(514, 61) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>0 Ti4>0 Ti5>0 Ti6>1 Ti7>1 Ri0>0 To0<0 To1<0 To2<0 Lo0<0 Bo0<1 Bo1<0 ]
  tran g24(.Z(w37), .I(B[15:12]));   //: @(266,85) /sn:0 /R:1 /w:[ 1 1 2 ] /ss:1
  tran g18(.Z(w29), .I(A[11:8]));   //: @(356,41) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: joint g10 (Cin) @(828, 206) /w:[ 2 -1 4 1 ]
  //: output g25 (GG) @(256,429) /sn:0 /w:[ 0 ]
  led g6 (.I(w32));   //: @(318,143) /sn:0 /w:[ 1 ] /type:0
  led g7 (.I(w9));   //: @(511,146) /sn:0 /w:[ 0 ] /type:0
  //: input g9 (Cin) @(900,206) /sn:0 /R:2 /w:[ 3 ]
  tran g22(.Z(w23), .I(B[7:4]));   //: @(611,84) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  //: input g12 (A) @(150,43) /sn:0 /w:[ 0 ]
  led g5 (.I(w39));   //: @(170,161) /sn:0 /w:[ 1 ] /type:0
  //: output g11 (Cout) @(153,345) /sn:0 /R:2 /w:[ 5 ]
  //: joint g14 (Cout) @(184, 346) /w:[ 1 -1 2 4 ]
  tran g19(.Z(w22), .I(A[7:4]));   //: @(553,41) /sn:0 /R:1 /w:[ 1 5 6 ] /ss:1
  tran g21(.Z(w1), .I(B[3:0]));   //: @(777,85) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  tran g20(.Z(w0), .I(A[3:0]));   //: @(719,41) /sn:0 /R:1 /w:[ 1 7 8 ] /ss:1
  CLA4 g0 (.B(w1), .A(w0), .Cin(Cin), .Cout(w10), .GG(w14), .PG(w13), .S(w2));   //: @(701, 157) /sz:(108, 57) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>5 Lo0<1 Bo0<1 Bo1<1 Bo2<1 ]
  concat g15 (.I0(w2), .I1(w3), .I2(w8), .I3(w15), .Z(S));   //: @(867,418) /sn:0 /w:[ 0 0 0 0 1 ] /dr:0
  //: input g13 (B) @(151,87) /sn:0 /w:[ 0 ]

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 {0}(461,53)(461,127)(354,127)(354,137){1}
wire w7;    //: /sn:0 {0}(454,193)(454,182)(393,182){1}
wire w4;    //: /sn:0 {0}(371,282)(371,233)(355,233)(355,223){1}
wire [15:0] w3;    //: /sn:0 {0}(120,283)(120,293)(316,293)(316,223){1}
wire w8;    //: /sn:0 {0}(416,281)(416,233)(376,233)(376,223){1}
wire [15:0] w2;    //: /sn:0 {0}(194,84)(194,127)(282,127)(282,137){1}
wire w5;    //: /sn:0 {0}(105,157)(105,177)(250,177){1}
//: enddecls

  led g4 (.I(w5));   //: @(105,150) /sn:0 /w:[ 0 ] /type:0
  led g3 (.I(w8));   //: @(416,288) /sn:0 /R:2 /w:[ 0 ] /type:0
  led g2 (.I(w4));   //: @(371,289) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: switch g1 (w7) @(454,207) /sn:0 /R:1 /w:[ 0 ] /st:1
  //: dip g6 (w2) @(194,74) /sn:0 /w:[ 0 ] /st:65535
  //: dip g7 (w6) @(461,43) /sn:0 /w:[ 0 ] /st:65535
  led g5 (.I(w3));   //: @(120,276) /sn:0 /w:[ 0 ] /type:2
  CLA16 g0 (.B(w6), .A(w2), .Cin(w7), .Cout(w5), .GG(w8), .PG(w4), .S(w3));   //: @(251, 138) /sz:(141, 84) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 Bo1<1 Bo2<1 ]

endmodule
