//: version "1.8.7"

module FA_alt(S, Co, B, A, Ci);
//: interface  /sz:(40, 40) /bd:[ Li0>A(12/40) Li1>B(26/40) Bi0>Ci(15/40) Ro0<S(22/40) Ro1<Co(31/40) ]
input B;    //: /sn:0 {0}(133,52)(133,126)(223,126){1}
//: {2}(227,126)(236,126){3}
//: {4}(225,128)(225,200)(232,200){5}
//: {6}(236,200)(251,200){7}
//: {8}(234,202)(234,221)(251,221){9}
input A;    //: /sn:0 {0}(115,52)(115,131)(204,131){1}
//: {2}(208,131)(236,131){3}
//: {4}(206,133)(206,205)(215,205){5}
//: {6}(219,205)(251,205){7}
//: {8}(217,207)(217,242)(251,242){9}
output Co;    //: /sn:0 {0}(352,224)(327,224){1}
input Ci;    //: /sn:0 {0}(251,226)(170,226)(170,161){1}
//: {2}(172,159)(308,159){3}
//: {4}(168,159)(123,159){5}
//: {6}(119,159)(98,159)(98,52){7}
//: {8}(121,161)(121,247)(251,247){9}
output S;    //: /sn:0 {0}(352,157)(329,157){1}
wire w16;    //: /sn:0 /dp:1 {0}(306,224)(272,224){1}
wire w3;    //: /sn:0 /dp:1 {0}(308,154)(267,154)(267,129)(257,129){1}
wire w18;    //: /sn:0 {0}(306,229)(282,229)(282,245)(272,245){1}
wire w8;    //: /sn:0 {0}(272,203)(296,203)(296,219)(306,219){1}
//: enddecls

  //: output g8 (S) @(349,157) /sn:0 /w:[ 0 ]
  and g4 (.I0(B), .I1(A), .Z(w8));   //: @(262,203) /sn:0 /delay:" 4" /w:[ 7 7 0 ]
  //: joint g16 (A) @(217, 205) /w:[ 6 -1 5 8 ]
  //: output g3 (Co) @(349,224) /sn:0 /w:[ 0 ]
  //: joint g17 (Ci) @(121, 159) /w:[ 5 -1 6 8 ]
  //: joint g2 (Ci) @(170, 159) /w:[ 2 -1 4 1 ]
  xnor g1 (.I0(w3), .I1(!Ci), .Z(S));   //: @(319,157) /sn:0 /delay:" 5" /w:[ 0 3 1 ]
  //: input g10 (B) @(133,50) /sn:0 /R:3 /w:[ 0 ]
  and g6 (.I0(A), .I1(Ci), .Z(w18));   //: @(262,245) /sn:0 /delay:" 4" /w:[ 9 9 1 ]
  //: input g9 (A) @(115,50) /sn:0 /R:3 /w:[ 0 ]
  or g7 (.I0(w8), .I1(w16), .I2(w18), .Z(Co));   //: @(317,224) /sn:0 /anc:1 /delay:" 4" /w:[ 1 0 0 1 ]
  //: joint g12 (B) @(225, 126) /w:[ 2 -1 1 4 ]
  //: joint g14 (B) @(234, 200) /w:[ 6 -1 5 8 ]
  //: input g11 (Ci) @(98,50) /sn:0 /R:3 /w:[ 7 ]
  and g5 (.I0(B), .I1(Ci), .Z(w16));   //: @(262,224) /sn:0 /delay:" 4" /w:[ 9 0 1 ]
  xor g0 (.I0(B), .I1(A), .Z(w3));   //: @(247,129) /sn:0 /delay:" 5" /w:[ 3 3 1 ]
  //: joint g13 (A) @(206, 131) /w:[ 2 -1 1 4 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(343,185)(315,185)(315,155)(305,155){1}
wire w0;    //: /sn:0 {0}(148,181)(200,181)(200,150)(263,150){1}
wire w3;    //: /sn:0 {0}(152,129)(198,129)(198,136)(263,136){1}
wire w1;    //: /sn:0 {0}(220,222)(270,222)(270,175)(279,175)(279,165){1}
wire w5;    //: /sn:0 {0}(416,82)(315,82)(315,146)(305,146){1}
//: enddecls

  //: switch g4 (w0) @(131,181) /sn:0 /w:[ 0 ] /st:0
  //: switch g3 (w3) @(135,129) /sn:0 /w:[ 0 ] /st:0
  led g2 (.I(w4));   //: @(350,185) /sn:0 /R:3 /w:[ 0 ] /type:0
  led g1 (.I(w5));   //: @(423,82) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: switch g5 (w1) @(203,222) /sn:0 /w:[ 0 ] /st:0
  FA_alt g0 (.B(w0), .A(w3), .Ci(w1), .Co(w4), .S(w5));   //: @(264, 124) /sz:(40, 40) /sn:0 /p:[ Li0>1 Li1>1 Bi0>1 Ro0<1 Ro1<1 ]

endmodule
