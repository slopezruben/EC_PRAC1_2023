//: version "1.8.7"

module PFA(Si, Gi, Ci, b, Pi, a);
//: interface  /sz:(100, 59) /bd:[ Ti0>b(61/100) Ti1>a(29/100) Ri0>Ci(28/59) Bo0<Pi(20/100) Bo1<Gi(52/100) Bo2<Si(83/100) ]
input b;    //: /sn:0 {0}(90,69)(103,69){1}
//: {2}(107,69)(155,69)(155,61)(159,61){3}
//: {4}(105,71)(105,104){5}
//: {6}(107,106)(243,106){7}
//: {8}(105,108)(105,136)(234,136){9}
output Gi;    //: /sn:0 /dp:1 {0}(255,134)(286,134){1}
output Si;    //: /sn:0 /dp:1 {0}(256,80)(283,80){1}
output Pi;    //: /sn:0 /dp:1 {0}(264,104)(288,104){1}
input Ci;    //: /sn:0 {0}(87,88)(225,88)(225,82)(235,82){1}
input a;    //: /sn:0 {0}(88,54)(116,54){1}
//: {2}(120,54)(151,54)(151,56)(159,56){3}
//: {4}(118,56)(118,99){5}
//: {6}(120,101)(243,101){7}
//: {8}(118,103)(118,131)(234,131){9}
wire w2;    //: /sn:0 {0}(180,59)(225,59)(225,77)(235,77){1}
//: enddecls

  //: output g4 (Si) @(280,80) /sn:0 /w:[ 1 ]
  or g8 (.I0(a), .I1(b), .Z(Pi));   //: @(254,104) /sn:0 /delay:" 4" /w:[ 7 7 0 ]
  //: output g3 (Gi) @(283,134) /sn:0 /w:[ 1 ]
  //: input g2 (Ci) @(85,88) /sn:0 /w:[ 0 ]
  //: input g1 (b) @(88,69) /sn:0 /w:[ 0 ]
  //: joint g10 (a) @(118, 54) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(a), .I1(b), .Z(w2));   //: @(170,59) /sn:0 /delay:" 5" /w:[ 3 3 0 ]
  xor g7 (.I0(w2), .I1(Ci), .Z(Si));   //: @(246,80) /sn:0 /delay:" 5" /w:[ 1 1 0 ]
  and g9 (.I0(a), .I1(b), .Z(Gi));   //: @(245,134) /sn:0 /delay:" 4" /w:[ 9 9 0 ]
  //: joint g12 (a) @(118, 101) /w:[ 6 5 -1 8 ]
  //: joint g11 (b) @(105, 69) /w:[ 2 -1 1 4 ]
  //: output g5 (Pi) @(285,104) /sn:0 /w:[ 1 ]
  //: input g0 (a) @(86,54) /sn:0 /w:[ 0 ]
  //: joint g13 (b) @(105, 106) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(215,91)(228,91)(228,142){1}
wire w7;    //: /sn:0 {0}(250,45)(260,45)(260,142){1}
wire w10;    //: /sn:0 {0}(251,242)(251,203){1}
wire w11;    //: /sn:0 {0}(219,242)(219,203){1}
wire w2;    //: /sn:0 /dp:1 {0}(300,171)(329,171)(329,189){1}
wire w9;    //: /sn:0 {0}(282,283)(282,203){1}
//: enddecls

  led g4 (.I(w9));   //: @(282,290) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: switch g3 (w2) @(329,203) /sn:0 /R:1 /w:[ 1 ] /st:0
  //: switch g2 (w7) @(233,45) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w6) @(198,91) /sn:0 /w:[ 0 ] /st:0
  led g6 (.I(w11));   //: @(219,249) /sn:0 /R:2 /w:[ 0 ] /type:0
  led g5 (.I(w10));   //: @(251,249) /sn:0 /R:2 /w:[ 0 ] /type:0
  PFA g0 (.b(w7), .a(w6), .Ci(w2), .Pi(w11), .Gi(w10), .Si(w9));   //: @(199, 143) /sz:(100, 59) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<1 Bo1<1 Bo2<1 ]

endmodule
