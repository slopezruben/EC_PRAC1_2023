//: version "1.8.7"

module main;    //: root_module
wire w6;    //: /sn:0 {0}(567,155)(530,155){1}
wire w7;    //: /sn:0 {0}(511,97)(511,137){1}
wire w8;    //: /sn:0 {0}(486,69)(486,137){1}
wire w5;    //: /sn:0 {0}(440,161)(469,161){1}
wire w9;    //: /sn:0 {0}(495,201)(495,179){1}
//: enddecls

  led g4 (.I(w5));   //: @(433,161) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: switch g3 (w6) @(585,155) /sn:0 /R:2 /w:[ 0 ] /st:1
  //: switch g2 (w7) @(511,84) /sn:0 /R:3 /w:[ 0 ] /st:1
  //: switch g1 (w8) @(486,56) /sn:0 /R:3 /w:[ 0 ] /st:1
  FA g7 (.B(w7), .A(w8), .Cin(w6), .Cout(w5), .S(w9));   //: @(470, 138) /sz:(59, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  led g5 (.I(w9));   //: @(495,208) /sn:0 /R:2 /w:[ 0 ] /type:0

endmodule

module FA(Cout, S, Cin, B, A);
//: interface  /sz:(59, 40) /bd:[ Ti0>A(16/59) Ti1>B(41/59) Ri0>Cin(17/40) Lo0<Cout(23/40) Bo0<S(25/59) ]
input B;    //: /sn:0 {0}(249,96)(296,96)(296,126){1}
input A;    //: /sn:0 {0}(193,113)(276,113)(276,126){1}
input Cin;    //: /sn:0 {0}(345,185)(345,76)(288,76){1}
output Cout;    //: /sn:0 {0}(323,329)(224,329)(224,286){1}
output S;    //: /sn:0 /dp:1 {0}(334,227)(334,264)(350,264){1}
wire w3;    //: /sn:0 /dp:1 {0}(222,265)(222,157)(267,157){1}
wire w0;    //: /sn:0 /dp:1 {0}(227,265)(227,255)(251,255)(251,216)(316,216){1}
wire w1;    //: /sn:0 {0}(325,185)(325,180)(285,180)(285,168){1}
//: enddecls

  //: output g4 (Cout) @(320,329) /sn:0 /w:[ 0 ]
  //: output g3 (S) @(347,264) /sn:0 /w:[ 1 ]
  //: input g2 (Cin) @(286,76) /sn:0 /w:[ 1 ]
  //: input g1 (B) @(247,96) /sn:0 /w:[ 0 ]
  HA g6 (.A(w1), .B(Cin), .C(w0), .S(S));   //: @(317, 186) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<1 Bo0<0 ]
  or g7 (.I0(w0), .I1(w3), .Z(Cout));   //: @(224,276) /sn:0 /R:3 /delay:" 4" /w:[ 0 0 1 ]
  HA g5 (.A(A), .B(B), .C(w3), .S(w1));   //: @(268, 127) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]
  //: input g0 (A) @(191,113) /sn:0 /w:[ 0 ]

endmodule
