//: version "1.8.7"

module RCA_4bits(Z, B, A);
//: interface  /sz:(111, 41) /bd:[ Ti0>A[3:0](41/111) Ti1>B[3:0](80/111) Bo0<Z[7:0](41/111) ]
input [3:0] B;    //: /sn:0 {0}(357,128)(373,128){1}
//: {2}(374,128)(568,128)(568,126)(618,126){3}
//: {4}(619,126)(713,126){5}
//: {6}(714,126)(789,126)(789,128)(798,128){7}
//: {8}(799,128)(876,128){9}
input [3:0] A;    //: /sn:0 {0}(378,82)(542,82){1}
//: {2}(543,82)(659,82){3}
//: {4}(660,82)(753,82){5}
//: {6}(754,82)(793,82){7}
//: {8}(794,82)(915,82)(915,72){9}
output [7:0] Z;    //: /sn:0 {0}(996,1089)(971,1089)(971,878)(961,878){1}
wire w16;    //: /sn:0 {0}(758,191)(758,330){1}
wire w13;    //: /sn:0 {0}(747,372)(747,903)(955,903){1}
wire w50;    //: /sn:0 {0}(33,677)(-47,677)(-47,679)(-57,679){1}
wire w34;    //: /sn:0 {0}(398,427)(398,476)(401,476)(401,486){1}
wire w39;    //: /sn:0 {0}(369,615)(369,624)(380,624)(380,634){1}
wire w3;    //: /sn:0 {0}(247,486)(247,429)(240,429)(240,419){1}
wire w36;    //: /sn:0 {0}(384,510)(301,510)(301,504)(291,504){1}
wire w22;    //: /sn:0 {0}(590,243)(590,327)(596,327)(596,337){1}
wire w0;    //: /sn:0 {0}(660,86)(660,104)(661,104)(661,110){1}
//: {2}(659,112)(454,112){3}
//: {4}(450,112)(237,112)(237,116){5}
//: {6}(235,118)(27,118)(27,586){7}
//: {8}(237,120)(237,398){9}
//: {10}(452,114)(452,271){11}
//: {12}(661,114)(661,175){13}
wire w20;    //: /sn:0 {0}(714,130)(714,208){1}
//: {2}(712,210)(594,210){3}
//: {4}(590,210)(463,210){5}
//: {6}(461,208)(461,191)(294,191)(294,252){7}
//: {8}(459,210)(457,210)(457,271){9}
//: {10}(592,212)(592,222){11}
//: {12}(714,212)(714,275){13}
wire w30;    //: /sn:0 {0}(599,468)(599,452)(563,452)(563,442){1}
wire w29;    //: /sn:0 {0}(301,384)(301,476)(272,476)(272,486){1}
wire w42;    //: /sn:0 {0}(52,517)(-76,517)(-76,661){1}
wire w37;    //: /sn:0 {0}(410,528)(410,624)(400,624)(400,634){1}
wire w18;    //: /sn:0 {0}(619,130)(619,136)(565,136)(565,297){1}
//: {2}(563,299)(402,299){3}
//: {4}(398,299)(341,299){5}
//: {6}(337,299)(153,299)(153,391){7}
//: {8}(339,301)(339,322)(242,322)(242,398){9}
//: {10}(400,301)(400,406){11}
//: {12}(565,301)(565,421){13}
wire w19;    //: /sn:0 {0}(478,269)(478,324)(471,324)(471,334){1}
wire w12;    //: /sn:0 {0}(729,361)(650,361)(650,355)(640,355){1}
wire w23;    //: /sn:0 {0}(455,292)(455,324)(446,324)(446,334){1}
wire w10;    //: /sn:0 {0}(796,192)(796,913)(955,913){1}
wire w54;    //: /sn:0 {0}(-92,703)(-92,853)(955,853){1}
wire w24;    //: /sn:0 {0}(579,361)(500,361)(500,352)(490,352){1}
wire w1;    //: /sn:0 {0}(619,468)(619,389)(605,389)(605,379){1}
wire w31;    //: /sn:0 {0}(292,273)(292,342){1}
wire w32;    //: /sn:0 {0}(590,499)(455,499)(455,504)(445,504){1}
wire w53;    //: /sn:0 {0}(-118,685)(-128,685)(-128,843)(955,843){1}
wire w46;    //: /sn:0 {0}(371,665)(270,665){1}
wire w52;    //: /sn:0 {0}(30,607)(30,643)(50,643)(50,653){1}
wire w27;    //: /sn:0 {0}(429,358)(327,358)(327,332)(312,332)(312,342){1}
wire w17;    //: /sn:0 {0}(664,196)(664,327)(621,327)(621,337){1}
wire w35;    //: /sn:0 {0}(374,132)(374,556)(384,556)(384,562){1}
//: {2}(382,564)(215,564){3}
//: {4}(211,564)(203,564)(203,600){5}
//: {6}(213,566)(213,576)(34,576){7}
//: {8}(30,576)(-113,576)(-113,594){9}
//: {10}(32,578)(32,586){11}
//: {12}(384,566)(384,577)(371,577)(371,594){13}
wire w33;    //: /sn:0 {0}(608,510)(608,893)(955,893){1}
wire w28;    //: /sn:0 {0}(455,376)(455,476)(426,476)(426,486){1}
wire w49;    //: /sn:0 {0}(201,621)(201,637)(226,637)(226,647){1}
wire w45;    //: /sn:0 {0}(209,671)(94,671){1}
wire w14;    //: /sn:0 {0}(754,86)(754,100)(755,100)(755,111){1}
//: {2}(753,113)(743,113)(743,120)(589,120){3}
//: {4}(585,120)(395,120)(395,169){5}
//: {6}(393,171)(198,171)(198,600){7}
//: {8}(395,173)(395,406){9}
//: {10}(587,122)(587,222){11}
//: {12}(755,115)(755,170){13}
wire w48;    //: /sn:0 {0}(235,689)(235,873)(955,873){1}
wire w41;    //: /sn:0 {0}(256,528)(256,637)(251,637)(251,647){1}
wire w11;    //: /sn:0 {0}(738,330)(738,306)(712,306)(712,296){1}
wire w2;    //: /sn:0 {0}(560,421)(560,397){1}
//: {2}(560,393)(560,98)(707,98){3}
//: {4}(711,98)(792,98){5}
//: {6}(794,96)(794,86){7}
//: {8}(794,100)(794,115)(793,115)(793,171){9}
//: {10}(709,100)(709,275){11}
//: {12}(558,395)(366,395)(366,594){13}
wire w47;    //: /sn:0 {0}(389,676)(389,883)(955,883){1}
wire w15;    //: /sn:0 {0}(543,86)(543,98){1}
//: {2}(541,100)(322,100){3}
//: {4}(318,100)(148,100)(148,224){5}
//: {6}(146,226)(-118,226)(-118,594){7}
//: {8}(148,228)(148,391){9}
//: {10}(320,102)(320,163)(289,163)(289,252){11}
//: {12}(543,102)(543,139)(475,139)(475,248){13}
wire w38;    //: /sn:0 {0}(151,412)(151,453)(63,453)(63,473)(69,473)(69,493){1}
wire w43;    //: /sn:0 {0}(78,535)(78,643)(75,643)(75,653){1}
wire w26;    //: /sn:0 {0}(283,373)(94,373)(94,493){1}
wire w9;    //: /sn:0 {0}(799,132)(799,134)(798,134)(798,142){1}
//: {2}(796,144)(762,144){3}
//: {4}(758,144)(668,144){5}
//: {6}(664,144)(480,144)(480,248){7}
//: {8}(666,146)(666,175){9}
//: {10}(760,146)(760,170){11}
//: {12}(798,146)(798,171){13}
wire w57;    //: /sn:0 {0}(-115,615)(-115,651)(-101,651)(-101,661){1}
wire w51;    //: /sn:0 {0}(59,695)(59,863)(955,863){1}
wire w40;    //: /sn:0 {0}(230,510)(123,510)(123,511)(113,511){1}
//: enddecls

  //: joint g75 (w35) @(213, 564) /w:[ 3 -1 4 6 ]
  HA g44 (.A(w31), .B(w27), .C(w26), .S(w29));   //: @(284, 343) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  HA g8 (.A(w11), .B(w16), .C(w12), .S(w13));   //: @(730, 331) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>1 Lo0<0 Bo0<0 ]
  and g4 (.I0(w2), .I1(w9), .Z(w10));   //: @(796,182) /sn:0 /R:3 /anc:1 /delay:" 4" /w:[ 9 13 0 ]
  //: joint g47 (w15) @(543, 100) /w:[ -1 1 2 12 ]
  //: comment g16 /dolink:0 /link:"" @(482,229) /sn:0 /R:3
  //: /line:"a3 * b0"
  //: /end
  concat g3 (.I0(w10), .I1(w13), .I2(w33), .I3(w47), .I4(w48), .I5(w51), .I6(w54), .I7(w53), .Z(Z));   //: @(960,878) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:0
  //: comment g26 /dolink:0 /link:"" @(-132,545) /sn:0 /R:3
  //: /line:"a3 * b3"
  //: /end
  //: comment g17 /dolink:0 /link:"" @(693,285) /sn:0 /R:3
  //: /line:"a0 * b1"
  //: /end
  //: output g2 (Z) @(993,1089) /sn:0 /w:[ 0 ]
  //: joint g74 (w0) @(237, 118) /w:[ -1 5 6 8 ]
  and g30 (.I0(w15), .I1(w9), .Z(w19));   //: @(478,259) /sn:0 /R:3 /delay:" 4" /w:[ 13 7 0 ]
  //: comment g23 /dolink:0 /link:"" @(351,597) /sn:0 /R:3
  //: /line:"a0 * b3"
  //: /end
  and g77 (.I0(w15), .I1(w35), .Z(w57));   //: @(-115,605) /sn:0 /R:3 /delay:" 4" /w:[ 7 9 0 ]
  FA g39 (.B(w17), .A(w22), .Cin(w12), .Cout(w24), .S(w1));   //: @(580, 338) /sz:(59, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  //: comment g24 /dolink:0 /link:"" @(150,596) /sn:0 /R:3
  //: /line:"a1 * b3"
  //: /end
  //: input g1 (B) @(355,128) /sn:0 /w:[ 0 ]
  //: joint g60 (w18) @(339, 299) /w:[ 5 -1 6 8 ]
  tran g29(.Z(w0), .I(A[2]));   //: @(660,80) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  HA g51 (.A(w30), .B(w1), .C(w32), .S(w33));   //: @(591, 469) /sz:(40, 40) /sn:0 /p:[ Ti0>0 Ti1>0 Lo0<0 Bo0<0 ]
  //: joint g70 (w14) @(395, 171) /w:[ -1 5 6 8 ]
  //: comment g18 /dolink:0 /link:"" @(262,279) /sn:0 /R:3
  //: /line:"a3 * b1"
  //: /end
  HA g65 (.A(w39), .B(w37), .C(w46), .S(w47));   //: @(372, 635) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<0 Bo0<0 ]
  //: comment g25 /dolink:0 /link:"" @(12,593) /sn:0 /R:3
  //: /line:"a2 * b3"
  //: /end
  //: comment g10 /dolink:0 /link:"" @(566,244) /sn:0 /R:3
  //: /line:"a1 * b1"
  //: /end
  and g64 (.I0(w2), .I1(w35), .Z(w39));   //: @(369,605) /sn:0 /R:3 /delay:" 4" /w:[ 13 13 0 ]
  FA g72 (.B(w43), .A(w52), .Cin(w45), .Cout(w50), .S(w51));   //: @(34, 654) /sz:(59, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g49 (w14) @(755, 113) /w:[ -1 1 2 12 ]
  tran g50(.Z(w18), .I(B[2]));   //: @(619,124) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g6(.Z(w2), .I(A[0]));   //: @(794,80) /sn:0 /R:1 /w:[ 7 7 8 ] /ss:1
  and g73 (.I0(w0), .I1(w35), .Z(w52));   //: @(30,597) /sn:0 /R:3 /delay:" 4" /w:[ 7 11 0 ]
  FA g68 (.B(w41), .A(w49), .Cin(w46), .Cout(w45), .S(w48));   //: @(210, 648) /sz:(59, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g58 (w18) @(400, 299) /w:[ 3 -1 4 10 ]
  and g56 (.I0(w0), .I1(w18), .Z(w3));   //: @(240,409) /sn:0 /R:3 /delay:" 4" /w:[ 9 9 1 ]
  tran g35(.Z(w20), .I(B[1]));   //: @(714,124) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  and g9 (.I0(w14), .I1(w9), .Z(w16));   //: @(758,181) /sn:0 /R:3 /delay:" 4" /w:[ 13 11 0 ]
  //: comment g7 /dolink:0 /link:"" @(812,171) /sn:0 /R:3
  //: /line:"a0 * b0"
  //: /end
  //: joint g71 (w35) @(384, 564) /w:[ -1 1 2 12 ]
  and g59 (.I0(w15), .I1(w18), .Z(w38));   //: @(151,402) /sn:0 /R:3 /delay:" 4" /w:[ 9 7 0 ]
  //: joint g31 (w9) @(666, 144) /w:[ 5 -1 6 8 ]
  //: comment g22 /dolink:0 /link:"" @(219,401) /sn:0 /R:3
  //: /line:"a2 * b2"
  //: /end
  tran g67(.Z(w35), .I(B[3]));   //: @(374,126) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g54 (w18) @(565, 299) /w:[ -1 1 2 12 ]
  and g45 (.I0(w15), .I1(w20), .Z(w31));   //: @(292,263) /sn:0 /R:3 /delay:" 4" /w:[ 11 7 0 ]
  //: joint g41 (w0) @(661, 112) /w:[ -1 1 2 12 ]
  and g36 (.I0(w14), .I1(w20), .Z(w22));   //: @(590,233) /sn:0 /R:3 /delay:" 4" /w:[ 11 11 0 ]
  and g33 (.I0(w2), .I1(w20), .Z(w11));   //: @(712,286) /sn:0 /R:3 /delay:" 4" /w:[ 11 13 1 ]
  and g69 (.I0(w14), .I1(w35), .Z(w49));   //: @(201,611) /sn:0 /R:3 /delay:" 4" /w:[ 7 5 0 ]
  and g52 (.I0(w14), .I1(w18), .Z(w34));   //: @(398,417) /sn:0 /R:3 /delay:" 4" /w:[ 9 11 0 ]
  //: joint g42 (w20) @(592, 210) /w:[ 3 -1 4 10 ]
  and g40 (.I0(w0), .I1(w20), .Z(w23));   //: @(455,282) /sn:0 /R:3 /delay:" 4" /w:[ 11 9 0 ]
  //: joint g66 (w2) @(560, 395) /w:[ -1 2 12 1 ]
  //: joint g12 (w9) @(798, 144) /w:[ -1 1 2 12 ]
  //: joint g57 (w0) @(452, 112) /w:[ 3 -1 4 10 ]
  //: joint g46 (w20) @(461, 210) /w:[ 5 6 8 -1 ]
  //: joint g34 (w2) @(794, 98) /w:[ -1 6 5 8 ]
  //: comment g28 /dolink:0 /link:"" @(745,196) /sn:0 /R:3
  //: /line:"a1*b0"
  //: /end
  //: comment g14 /dolink:0 /link:"" @(385,259) /sn:0 /R:3
  //: /line:"a2 * b1"
  //: /end
  tran g11(.Z(w14), .I(A[1]));   //: @(754,80) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g5(.Z(w9), .I(B[0]));   //: @(799,126) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: joint g61 (w15) @(320, 100) /w:[ 3 -1 4 10 ]
  //: comment g21 /dolink:0 /link:"" @(104,345) /sn:0 /R:3
  //: /line:"a3*b2"
  //: /end
  //: comment g19 /dolink:0 /link:"" @(551,428) /sn:0 /R:3
  //: /line:"a0*b2"
  //: /line:""
  //: /end
  //: joint g79 (w15) @(148, 226) /w:[ -1 5 6 8 ]
  //: joint g78 (w35) @(32, 576) /w:[ 7 -1 8 10 ]
  tran g32(.Z(w15), .I(A[3]));   //: @(543,80) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: comment g20 /dolink:0 /link:"" @(382,425) /sn:0 /R:3
  //: /line:"a1 * b2"
  //: /end
  FA g63 (.B(w26), .A(w38), .Cin(w40), .Cout(w42), .S(w43));   //: @(53, 494) /sz:(59, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g43 (.B(w19), .A(w23), .Cin(w24), .Cout(w27), .S(w28));   //: @(430, 335) /sz:(59, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g38 (w20) @(714, 210) /w:[ -1 1 2 12 ]
  //: comment g15 /dolink:0 /link:"" @(648,192) /sn:0 /R:3
  //: /line:"a2 * b0"
  //: /end
  //: input g0 (A) @(376,82) /sn:0 /w:[ 0 ]
  and g48 (.I0(w2), .I1(w18), .Z(w30));   //: @(563,432) /sn:0 /R:3 /delay:" 4" /w:[ 0 13 1 ]
  //: joint g27 (w9) @(760, 144) /w:[ 3 -1 4 10 ]
  FA g62 (.B(w29), .A(w3), .Cin(w36), .Cout(w40), .S(w41));   //: @(231, 487) /sz:(59, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g37 (w2) @(709, 98) /w:[ 4 -1 3 10 ]
  FA g55 (.B(w28), .A(w34), .Cin(w32), .Cout(w36), .S(w37));   //: @(385, 487) /sz:(59, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g76 (.B(w42), .A(w57), .Cin(w50), .Cout(w53), .S(w54));   //: @(-117, 662) /sz:(59, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  //: joint g53 (w14) @(587, 120) /w:[ 3 -1 4 10 ]
  and g13 (.I0(w0), .I1(w9), .Z(w17));   //: @(664,186) /sn:0 /R:3 /delay:" 4" /w:[ 13 9 0 ]

endmodule

module main;    //: root_module
wire [3:0] w4;    //: /sn:0 {0}(315,50)(310,50)(310,137){1}
wire [7:0] w0;    //: /sn:0 {0}(352,261)(271,261)(271,180){1}
wire [3:0] w3;    //: /sn:0 {0}(165,39)(155,39)(155,54)(271,54)(271,137){1}
//: enddecls

  led g3 (.I(w0));   //: @(359,261) /sn:0 /R:3 /w:[ 0 ] /type:3
  //: dip g2 (w4) @(353,50) /sn:0 /R:3 /w:[ 0 ] /st:10
  //: dip g1 (w3) @(203,39) /sn:0 /R:3 /w:[ 0 ] /st:10
  RCA_4bits g0 (.B(w4), .A(w3), .Z(w0));   //: @(230, 138) /sz:(111, 41) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 ]

endmodule
